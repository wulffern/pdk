magic
tech sky130A
magscale 1 2
timestamp 1665766018
<< nwell >>
rect 0 0 816 240
<< pmos >>
rect 95 36 125 204
rect 181 36 211 204
rect 267 36 297 204
rect 353 36 383 204
rect 439 36 469 204
rect 525 36 555 204
rect 611 36 641 204
rect 697 36 727 204
<< pdiff >>
rect 42 173 95 204
rect 42 139 50 173
rect 84 139 95 173
rect 42 101 95 139
rect 42 67 50 101
rect 84 67 95 101
rect 42 36 95 67
rect 125 173 181 204
rect 125 139 136 173
rect 170 139 181 173
rect 125 101 181 139
rect 125 67 136 101
rect 170 67 181 101
rect 125 36 181 67
rect 211 173 267 204
rect 211 139 222 173
rect 256 139 267 173
rect 211 101 267 139
rect 211 67 222 101
rect 256 67 267 101
rect 211 36 267 67
rect 297 173 353 204
rect 297 139 308 173
rect 342 139 353 173
rect 297 101 353 139
rect 297 67 308 101
rect 342 67 353 101
rect 297 36 353 67
rect 383 173 439 204
rect 383 139 394 173
rect 428 139 439 173
rect 383 101 439 139
rect 383 67 394 101
rect 428 67 439 101
rect 383 36 439 67
rect 469 173 525 204
rect 469 139 480 173
rect 514 139 525 173
rect 469 101 525 139
rect 469 67 480 101
rect 514 67 525 101
rect 469 36 525 67
rect 555 173 611 204
rect 555 139 566 173
rect 600 139 611 173
rect 555 101 611 139
rect 555 67 566 101
rect 600 67 611 101
rect 555 36 611 67
rect 641 173 697 204
rect 641 139 652 173
rect 686 139 697 173
rect 641 101 697 139
rect 641 67 652 101
rect 686 67 697 101
rect 641 36 697 67
rect 727 173 780 204
rect 727 139 738 173
rect 772 139 780 173
rect 727 101 780 139
rect 727 67 738 101
rect 772 67 780 101
rect 727 36 780 67
<< pdiffc >>
rect 50 139 84 173
rect 50 67 84 101
rect 136 139 170 173
rect 136 67 170 101
rect 222 139 256 173
rect 222 67 256 101
rect 308 139 342 173
rect 308 67 342 101
rect 394 139 428 173
rect 394 67 428 101
rect 480 139 514 173
rect 480 67 514 101
rect 566 139 600 173
rect 566 67 600 101
rect 652 139 686 173
rect 652 67 686 101
rect 738 139 772 173
rect 738 67 772 101
<< poly >>
rect 95 287 727 303
rect 95 253 156 287
rect 190 253 224 287
rect 258 253 292 287
rect 326 253 360 287
rect 394 253 428 287
rect 462 253 496 287
rect 530 253 564 287
rect 598 253 632 287
rect 666 253 727 287
rect 95 230 727 253
rect 95 204 125 230
rect 181 204 211 230
rect 267 204 297 230
rect 353 204 383 230
rect 439 204 469 230
rect 525 204 555 230
rect 611 204 641 230
rect 697 204 727 230
rect 95 10 125 36
rect 181 10 211 36
rect 267 10 297 36
rect 353 10 383 36
rect 439 10 469 36
rect 525 10 555 36
rect 611 10 641 36
rect 697 10 727 36
<< polycont >>
rect 156 253 190 287
rect 224 253 258 287
rect 292 253 326 287
rect 360 253 394 287
rect 428 253 462 287
rect 496 253 530 287
rect 564 253 598 287
rect 632 253 666 287
<< locali >>
rect 140 287 682 303
rect 140 253 142 287
rect 190 253 214 287
rect 258 253 286 287
rect 326 253 358 287
rect 394 253 428 287
rect 464 253 496 287
rect 536 253 564 287
rect 608 253 632 287
rect 680 253 682 287
rect 140 235 682 253
rect 50 173 84 189
rect 50 101 84 139
rect 50 51 84 67
rect 136 173 170 189
rect 136 101 170 139
rect 136 51 170 67
rect 222 173 256 189
rect 222 101 256 139
rect 222 51 256 67
rect 308 173 342 189
rect 308 101 342 139
rect 308 51 342 67
rect 394 173 428 189
rect 394 101 428 139
rect 394 51 428 67
rect 480 173 514 189
rect 480 101 514 139
rect 480 51 514 67
rect 566 173 600 189
rect 566 101 600 139
rect 566 51 600 67
rect 652 173 686 189
rect 652 101 686 139
rect 652 51 686 67
rect 738 173 772 189
rect 738 101 772 139
rect 738 51 772 67
<< viali >>
rect 142 253 156 287
rect 156 253 176 287
rect 214 253 224 287
rect 224 253 248 287
rect 286 253 292 287
rect 292 253 320 287
rect 358 253 360 287
rect 360 253 392 287
rect 430 253 462 287
rect 462 253 464 287
rect 502 253 530 287
rect 530 253 536 287
rect 574 253 598 287
rect 598 253 608 287
rect 646 253 666 287
rect 666 253 680 287
rect 50 139 84 173
rect 50 67 84 101
rect 136 139 170 173
rect 136 67 170 101
rect 222 139 256 173
rect 222 67 256 101
rect 308 139 342 173
rect 308 67 342 101
rect 394 139 428 173
rect 394 67 428 101
rect 480 139 514 173
rect 480 67 514 101
rect 566 139 600 173
rect 566 67 600 101
rect 652 139 686 173
rect 652 67 686 101
rect 738 139 772 173
rect 738 67 772 101
<< metal1 >>
rect 130 287 692 299
rect 130 253 142 287
rect 176 253 214 287
rect 248 253 286 287
rect 320 253 358 287
rect 392 253 430 287
rect 464 253 502 287
rect 536 253 574 287
rect 608 253 646 287
rect 680 253 692 287
rect 130 241 692 253
rect 44 173 90 189
rect 44 139 50 173
rect 84 139 90 173
rect 44 101 90 139
rect 44 67 50 101
rect 84 67 90 101
rect 44 -29 90 67
rect 127 178 179 189
rect 127 114 179 126
rect 127 51 179 62
rect 216 173 262 189
rect 216 139 222 173
rect 256 139 262 173
rect 216 101 262 139
rect 216 67 222 101
rect 256 67 262 101
rect 216 -29 262 67
rect 299 178 351 189
rect 299 114 351 126
rect 299 51 351 62
rect 388 173 434 189
rect 388 139 394 173
rect 428 139 434 173
rect 388 101 434 139
rect 388 67 394 101
rect 428 67 434 101
rect 388 -29 434 67
rect 471 178 523 189
rect 471 114 523 126
rect 471 51 523 62
rect 560 173 606 189
rect 560 139 566 173
rect 600 139 606 173
rect 560 101 606 139
rect 560 67 566 101
rect 600 67 606 101
rect 560 -29 606 67
rect 643 178 695 189
rect 643 114 695 126
rect 643 51 695 62
rect 732 173 778 189
rect 732 139 738 173
rect 772 139 778 173
rect 732 101 778 139
rect 732 67 738 101
rect 772 67 778 101
rect 732 -29 778 67
rect 44 -89 778 -29
<< via1 >>
rect 127 173 179 178
rect 127 139 136 173
rect 136 139 170 173
rect 170 139 179 173
rect 127 126 179 139
rect 127 101 179 114
rect 127 67 136 101
rect 136 67 170 101
rect 170 67 179 101
rect 127 62 179 67
rect 299 173 351 178
rect 299 139 308 173
rect 308 139 342 173
rect 342 139 351 173
rect 299 126 351 139
rect 299 101 351 114
rect 299 67 308 101
rect 308 67 342 101
rect 342 67 351 101
rect 299 62 351 67
rect 471 173 523 178
rect 471 139 480 173
rect 480 139 514 173
rect 514 139 523 173
rect 471 126 523 139
rect 471 101 523 114
rect 471 67 480 101
rect 480 67 514 101
rect 514 67 523 101
rect 471 62 523 67
rect 643 173 695 178
rect 643 139 652 173
rect 652 139 686 173
rect 686 139 695 173
rect 643 126 695 139
rect 643 101 695 114
rect 643 67 652 101
rect 652 67 686 101
rect 686 67 695 101
rect 643 62 695 67
<< metal2 >>
rect 120 188 186 197
rect 120 132 125 188
rect 181 132 186 188
rect 120 126 127 132
rect 179 126 186 132
rect 120 114 186 126
rect 120 108 127 114
rect 179 108 186 114
rect 120 52 125 108
rect 181 52 186 108
rect 120 43 186 52
rect 292 188 358 197
rect 292 132 297 188
rect 353 132 358 188
rect 292 126 299 132
rect 351 126 358 132
rect 292 114 358 126
rect 292 108 299 114
rect 351 108 358 114
rect 292 52 297 108
rect 353 52 358 108
rect 292 43 358 52
rect 464 188 530 197
rect 464 132 469 188
rect 525 132 530 188
rect 464 126 471 132
rect 523 126 530 132
rect 464 114 530 126
rect 464 108 471 114
rect 523 108 530 114
rect 464 52 469 108
rect 525 52 530 108
rect 464 43 530 52
rect 636 188 702 197
rect 636 132 641 188
rect 697 132 702 188
rect 636 126 643 132
rect 695 126 702 132
rect 636 114 702 126
rect 636 108 643 114
rect 695 108 702 114
rect 636 52 641 108
rect 697 52 702 108
rect 636 43 702 52
<< via2 >>
rect 125 178 181 188
rect 125 132 127 178
rect 127 132 179 178
rect 179 132 181 178
rect 125 62 127 108
rect 127 62 179 108
rect 179 62 181 108
rect 125 52 181 62
rect 297 178 353 188
rect 297 132 299 178
rect 299 132 351 178
rect 351 132 353 178
rect 297 62 299 108
rect 299 62 351 108
rect 351 62 353 108
rect 297 52 353 62
rect 469 178 525 188
rect 469 132 471 178
rect 471 132 523 178
rect 523 132 525 178
rect 469 62 471 108
rect 471 62 523 108
rect 523 62 525 108
rect 469 52 525 62
rect 641 178 697 188
rect 641 132 643 178
rect 643 132 695 178
rect 695 132 697 178
rect 641 62 643 108
rect 643 62 695 108
rect 695 62 697 108
rect 641 52 697 62
<< metal3 >>
rect 120 188 702 197
rect 120 132 125 188
rect 181 132 297 188
rect 353 132 469 188
rect 525 132 641 188
rect 697 132 702 188
rect 120 131 702 132
rect 120 108 186 131
rect 120 52 125 108
rect 181 52 186 108
rect 120 43 186 52
rect 292 108 358 131
rect 292 52 297 108
rect 353 52 358 108
rect 292 43 358 52
rect 464 108 530 131
rect 464 52 469 108
rect 525 52 530 108
rect 464 43 530 52
rect 636 108 702 131
rect 636 52 641 108
rect 697 52 702 108
rect 636 43 702 52
<< labels >>
flabel metal3 s 120 131 702 197 0 FreeSans 400 0 0 0 DRAIN
port 1 nsew
flabel metal1 s 44 -89 778 -29 0 FreeSans 400 0 0 0 SOURCE
port 2 nsew
flabel metal1 s 130 241 692 299 0 FreeSans 400 0 0 0 GATE
port 3 nsew
flabel nwell s 85 232 91 237 0 FreeSans 400 0 0 0 BULK
port 4 nsew
<< properties >>
string GDS_END 9221966
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9210038
string path 1.675 4.725 1.675 -2.225 
<< end >>
