/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/parameters/slow_70p.spice