magic
tech sky130A
magscale 1 2
timestamp 1665766018
<< nwell >>
rect 0 0 826 980
<< pmos >>
rect 171 189 201 791
rect 257 189 293 791
rect 349 189 385 791
rect 441 189 477 791
rect 533 189 569 791
rect 625 189 655 791
<< pdiff >>
rect 111 779 171 791
rect 111 745 126 779
rect 160 745 171 779
rect 111 711 171 745
rect 111 677 126 711
rect 160 677 171 711
rect 111 643 171 677
rect 111 609 126 643
rect 160 609 171 643
rect 111 575 171 609
rect 111 541 126 575
rect 160 541 171 575
rect 111 507 171 541
rect 111 473 126 507
rect 160 473 171 507
rect 111 439 171 473
rect 111 405 126 439
rect 160 405 171 439
rect 111 371 171 405
rect 111 337 126 371
rect 160 337 171 371
rect 111 303 171 337
rect 111 269 126 303
rect 160 269 171 303
rect 111 235 171 269
rect 111 201 126 235
rect 160 201 171 235
rect 111 189 171 201
rect 201 779 257 791
rect 201 745 212 779
rect 246 745 257 779
rect 201 711 257 745
rect 201 677 212 711
rect 246 677 257 711
rect 201 643 257 677
rect 201 609 212 643
rect 246 609 257 643
rect 201 575 257 609
rect 201 541 212 575
rect 246 541 257 575
rect 201 507 257 541
rect 201 473 212 507
rect 246 473 257 507
rect 201 439 257 473
rect 201 405 212 439
rect 246 405 257 439
rect 201 371 257 405
rect 201 337 212 371
rect 246 337 257 371
rect 201 303 257 337
rect 201 269 212 303
rect 246 269 257 303
rect 201 235 257 269
rect 201 201 212 235
rect 246 201 257 235
rect 201 189 257 201
rect 293 779 349 791
rect 293 745 304 779
rect 338 745 349 779
rect 293 711 349 745
rect 293 677 304 711
rect 338 677 349 711
rect 293 643 349 677
rect 293 609 304 643
rect 338 609 349 643
rect 293 575 349 609
rect 293 541 304 575
rect 338 541 349 575
rect 293 507 349 541
rect 293 473 304 507
rect 338 473 349 507
rect 293 439 349 473
rect 293 405 304 439
rect 338 405 349 439
rect 293 371 349 405
rect 293 337 304 371
rect 338 337 349 371
rect 293 303 349 337
rect 293 269 304 303
rect 338 269 349 303
rect 293 235 349 269
rect 293 201 304 235
rect 338 201 349 235
rect 293 189 349 201
rect 385 779 441 791
rect 385 745 396 779
rect 430 745 441 779
rect 385 711 441 745
rect 385 677 396 711
rect 430 677 441 711
rect 385 643 441 677
rect 385 609 396 643
rect 430 609 441 643
rect 385 575 441 609
rect 385 541 396 575
rect 430 541 441 575
rect 385 507 441 541
rect 385 473 396 507
rect 430 473 441 507
rect 385 439 441 473
rect 385 405 396 439
rect 430 405 441 439
rect 385 371 441 405
rect 385 337 396 371
rect 430 337 441 371
rect 385 303 441 337
rect 385 269 396 303
rect 430 269 441 303
rect 385 235 441 269
rect 385 201 396 235
rect 430 201 441 235
rect 385 189 441 201
rect 477 779 533 791
rect 477 745 488 779
rect 522 745 533 779
rect 477 711 533 745
rect 477 677 488 711
rect 522 677 533 711
rect 477 643 533 677
rect 477 609 488 643
rect 522 609 533 643
rect 477 575 533 609
rect 477 541 488 575
rect 522 541 533 575
rect 477 507 533 541
rect 477 473 488 507
rect 522 473 533 507
rect 477 439 533 473
rect 477 405 488 439
rect 522 405 533 439
rect 477 371 533 405
rect 477 337 488 371
rect 522 337 533 371
rect 477 303 533 337
rect 477 269 488 303
rect 522 269 533 303
rect 477 235 533 269
rect 477 201 488 235
rect 522 201 533 235
rect 477 189 533 201
rect 569 779 625 791
rect 569 745 580 779
rect 614 745 625 779
rect 569 711 625 745
rect 569 677 580 711
rect 614 677 625 711
rect 569 643 625 677
rect 569 609 580 643
rect 614 609 625 643
rect 569 575 625 609
rect 569 541 580 575
rect 614 541 625 575
rect 569 507 625 541
rect 569 473 580 507
rect 614 473 625 507
rect 569 439 625 473
rect 569 405 580 439
rect 614 405 625 439
rect 569 371 625 405
rect 569 337 580 371
rect 614 337 625 371
rect 569 303 625 337
rect 569 269 580 303
rect 614 269 625 303
rect 569 235 625 269
rect 569 201 580 235
rect 614 201 625 235
rect 569 189 625 201
rect 655 779 715 791
rect 655 745 666 779
rect 700 745 715 779
rect 655 711 715 745
rect 655 677 666 711
rect 700 677 715 711
rect 655 643 715 677
rect 655 609 666 643
rect 700 609 715 643
rect 655 575 715 609
rect 655 541 666 575
rect 700 541 715 575
rect 655 507 715 541
rect 655 473 666 507
rect 700 473 715 507
rect 655 439 715 473
rect 655 405 666 439
rect 700 405 715 439
rect 655 371 715 405
rect 655 337 666 371
rect 700 337 715 371
rect 655 303 715 337
rect 655 269 666 303
rect 700 269 715 303
rect 655 235 715 269
rect 655 201 666 235
rect 700 201 715 235
rect 655 189 715 201
<< pdiffc >>
rect 126 745 160 779
rect 126 677 160 711
rect 126 609 160 643
rect 126 541 160 575
rect 126 473 160 507
rect 126 405 160 439
rect 126 337 160 371
rect 126 269 160 303
rect 126 201 160 235
rect 212 745 246 779
rect 212 677 246 711
rect 212 609 246 643
rect 212 541 246 575
rect 212 473 246 507
rect 212 405 246 439
rect 212 337 246 371
rect 212 269 246 303
rect 212 201 246 235
rect 304 745 338 779
rect 304 677 338 711
rect 304 609 338 643
rect 304 541 338 575
rect 304 473 338 507
rect 304 405 338 439
rect 304 337 338 371
rect 304 269 338 303
rect 304 201 338 235
rect 396 745 430 779
rect 396 677 430 711
rect 396 609 430 643
rect 396 541 430 575
rect 396 473 430 507
rect 396 405 430 439
rect 396 337 430 371
rect 396 269 430 303
rect 396 201 430 235
rect 488 745 522 779
rect 488 677 522 711
rect 488 609 522 643
rect 488 541 522 575
rect 488 473 522 507
rect 488 405 522 439
rect 488 337 522 371
rect 488 269 522 303
rect 488 201 522 235
rect 580 745 614 779
rect 580 677 614 711
rect 580 609 614 643
rect 580 541 614 575
rect 580 473 614 507
rect 580 405 614 439
rect 580 337 614 371
rect 580 269 614 303
rect 580 201 614 235
rect 666 745 700 779
rect 666 677 700 711
rect 666 609 700 643
rect 666 541 700 575
rect 666 473 700 507
rect 666 405 700 439
rect 666 337 700 371
rect 666 269 700 303
rect 666 201 700 235
<< nsubdiff >>
rect 41 779 111 791
rect 41 745 58 779
rect 92 745 111 779
rect 41 711 111 745
rect 41 677 58 711
rect 92 677 111 711
rect 41 643 111 677
rect 41 609 58 643
rect 92 609 111 643
rect 41 575 111 609
rect 41 541 58 575
rect 92 541 111 575
rect 41 507 111 541
rect 41 473 58 507
rect 92 473 111 507
rect 41 439 111 473
rect 41 405 58 439
rect 92 405 111 439
rect 41 371 111 405
rect 41 337 58 371
rect 92 337 111 371
rect 41 303 111 337
rect 41 269 58 303
rect 92 269 111 303
rect 41 235 111 269
rect 41 201 58 235
rect 92 201 111 235
rect 41 189 111 201
rect 715 779 785 791
rect 715 745 734 779
rect 768 745 785 779
rect 715 711 785 745
rect 715 677 734 711
rect 768 677 785 711
rect 715 643 785 677
rect 715 609 734 643
rect 768 609 785 643
rect 715 575 785 609
rect 715 541 734 575
rect 768 541 785 575
rect 715 507 785 541
rect 715 473 734 507
rect 768 473 785 507
rect 715 439 785 473
rect 715 405 734 439
rect 768 405 785 439
rect 715 371 785 405
rect 715 337 734 371
rect 768 337 785 371
rect 715 303 785 337
rect 715 269 734 303
rect 768 269 785 303
rect 715 235 785 269
rect 715 201 734 235
rect 768 201 785 235
rect 715 189 785 201
<< nsubdiffcont >>
rect 58 745 92 779
rect 58 677 92 711
rect 58 609 92 643
rect 58 541 92 575
rect 58 473 92 507
rect 58 405 92 439
rect 58 337 92 371
rect 58 269 92 303
rect 58 201 92 235
rect 734 745 768 779
rect 734 677 768 711
rect 734 609 768 643
rect 734 541 768 575
rect 734 473 768 507
rect 734 405 768 439
rect 734 337 768 371
rect 734 269 768 303
rect 734 201 768 235
<< poly >>
rect 243 959 583 980
rect 116 873 201 889
rect 116 839 132 873
rect 166 839 201 873
rect 243 857 260 959
rect 566 857 583 959
rect 243 841 583 857
rect 625 873 710 889
rect 116 823 201 839
rect 171 791 201 823
rect 257 791 293 841
rect 349 791 385 841
rect 441 791 477 841
rect 533 791 569 841
rect 625 839 660 873
rect 694 839 710 873
rect 625 823 710 839
rect 625 791 655 823
rect 171 157 201 189
rect 116 141 201 157
rect 116 107 132 141
rect 166 107 201 141
rect 257 139 293 189
rect 349 139 385 189
rect 441 139 477 189
rect 533 139 569 189
rect 625 157 655 189
rect 625 141 710 157
rect 116 91 201 107
rect 243 123 583 139
rect 243 21 260 123
rect 566 21 583 123
rect 625 107 660 141
rect 694 107 710 141
rect 625 91 710 107
rect 243 0 583 21
<< polycont >>
rect 132 839 166 873
rect 260 857 566 959
rect 660 839 694 873
rect 132 107 166 141
rect 260 21 566 123
rect 660 107 694 141
<< locali >>
rect 238 961 588 980
rect 116 873 182 889
rect 116 839 132 873
rect 166 839 182 873
rect 238 855 252 961
rect 574 855 588 961
rect 238 841 588 855
rect 644 873 710 889
rect 116 823 182 839
rect 644 839 660 873
rect 694 839 710 873
rect 644 823 710 839
rect 116 795 160 823
rect 666 795 710 823
rect 41 779 160 795
rect 41 745 58 779
rect 92 759 126 779
rect 94 745 126 759
rect 41 725 60 745
rect 94 725 160 745
rect 41 711 160 725
rect 41 677 58 711
rect 92 687 126 711
rect 94 677 126 687
rect 41 653 60 677
rect 94 653 160 677
rect 41 643 160 653
rect 41 609 58 643
rect 92 615 126 643
rect 94 609 126 615
rect 41 581 60 609
rect 94 581 160 609
rect 41 575 160 581
rect 41 541 58 575
rect 92 543 126 575
rect 94 541 126 543
rect 41 509 60 541
rect 94 509 160 541
rect 41 507 160 509
rect 41 473 58 507
rect 92 473 126 507
rect 41 471 160 473
rect 41 439 60 471
rect 94 439 160 471
rect 41 405 58 439
rect 94 437 126 439
rect 92 405 126 437
rect 41 399 160 405
rect 41 371 60 399
rect 94 371 160 399
rect 41 337 58 371
rect 94 365 126 371
rect 92 337 126 365
rect 41 327 160 337
rect 41 303 60 327
rect 94 303 160 327
rect 41 269 58 303
rect 94 293 126 303
rect 92 269 126 293
rect 41 255 160 269
rect 41 235 60 255
rect 94 235 160 255
rect 41 201 58 235
rect 94 221 126 235
rect 92 201 126 221
rect 41 185 160 201
rect 212 779 246 795
rect 212 711 246 725
rect 212 643 246 653
rect 212 575 246 581
rect 212 507 246 509
rect 212 471 246 473
rect 212 399 246 405
rect 212 327 246 337
rect 212 255 246 269
rect 212 185 246 201
rect 304 779 338 795
rect 304 711 338 725
rect 304 643 338 653
rect 304 575 338 581
rect 304 507 338 509
rect 304 471 338 473
rect 304 399 338 405
rect 304 327 338 337
rect 304 255 338 269
rect 304 185 338 201
rect 396 779 430 795
rect 396 711 430 725
rect 396 643 430 653
rect 396 575 430 581
rect 396 507 430 509
rect 396 471 430 473
rect 396 399 430 405
rect 396 327 430 337
rect 396 255 430 269
rect 396 185 430 201
rect 488 779 522 795
rect 488 711 522 725
rect 488 643 522 653
rect 488 575 522 581
rect 488 507 522 509
rect 488 471 522 473
rect 488 399 522 405
rect 488 327 522 337
rect 488 255 522 269
rect 488 185 522 201
rect 580 779 614 795
rect 580 711 614 725
rect 580 643 614 653
rect 580 575 614 581
rect 580 507 614 509
rect 580 471 614 473
rect 580 399 614 405
rect 580 327 614 337
rect 580 255 614 269
rect 580 185 614 201
rect 666 779 785 795
rect 700 759 734 779
rect 700 745 732 759
rect 768 745 785 779
rect 666 725 732 745
rect 766 725 785 745
rect 666 711 785 725
rect 700 687 734 711
rect 700 677 732 687
rect 768 677 785 711
rect 666 653 732 677
rect 766 653 785 677
rect 666 643 785 653
rect 700 615 734 643
rect 700 609 732 615
rect 768 609 785 643
rect 666 581 732 609
rect 766 581 785 609
rect 666 575 785 581
rect 700 543 734 575
rect 700 541 732 543
rect 768 541 785 575
rect 666 509 732 541
rect 766 509 785 541
rect 666 507 785 509
rect 700 473 734 507
rect 768 473 785 507
rect 666 471 785 473
rect 666 439 732 471
rect 766 439 785 471
rect 700 437 732 439
rect 700 405 734 437
rect 768 405 785 439
rect 666 399 785 405
rect 666 371 732 399
rect 766 371 785 399
rect 700 365 732 371
rect 700 337 734 365
rect 768 337 785 371
rect 666 327 785 337
rect 666 303 732 327
rect 766 303 785 327
rect 700 293 732 303
rect 700 269 734 293
rect 768 269 785 303
rect 666 255 785 269
rect 666 235 732 255
rect 766 235 785 255
rect 700 221 732 235
rect 700 201 734 221
rect 768 201 785 235
rect 666 185 785 201
rect 116 157 160 185
rect 666 157 710 185
rect 116 141 182 157
rect 116 107 132 141
rect 166 107 182 141
rect 644 141 710 157
rect 116 91 182 107
rect 238 125 588 139
rect 238 19 252 125
rect 574 19 588 125
rect 644 107 660 141
rect 694 107 710 141
rect 644 91 710 107
rect 238 0 588 19
<< viali >>
rect 252 959 574 961
rect 252 857 260 959
rect 260 857 566 959
rect 566 857 574 959
rect 252 855 574 857
rect 60 745 92 759
rect 92 745 94 759
rect 60 725 94 745
rect 60 677 92 687
rect 92 677 94 687
rect 60 653 94 677
rect 60 609 92 615
rect 92 609 94 615
rect 60 581 94 609
rect 60 541 92 543
rect 92 541 94 543
rect 60 509 94 541
rect 60 439 94 471
rect 60 437 92 439
rect 92 437 94 439
rect 60 371 94 399
rect 60 365 92 371
rect 92 365 94 371
rect 60 303 94 327
rect 60 293 92 303
rect 92 293 94 303
rect 60 235 94 255
rect 60 221 92 235
rect 92 221 94 235
rect 212 745 246 759
rect 212 725 246 745
rect 212 677 246 687
rect 212 653 246 677
rect 212 609 246 615
rect 212 581 246 609
rect 212 541 246 543
rect 212 509 246 541
rect 212 439 246 471
rect 212 437 246 439
rect 212 371 246 399
rect 212 365 246 371
rect 212 303 246 327
rect 212 293 246 303
rect 212 235 246 255
rect 212 221 246 235
rect 304 745 338 759
rect 304 725 338 745
rect 304 677 338 687
rect 304 653 338 677
rect 304 609 338 615
rect 304 581 338 609
rect 304 541 338 543
rect 304 509 338 541
rect 304 439 338 471
rect 304 437 338 439
rect 304 371 338 399
rect 304 365 338 371
rect 304 303 338 327
rect 304 293 338 303
rect 304 235 338 255
rect 304 221 338 235
rect 396 745 430 759
rect 396 725 430 745
rect 396 677 430 687
rect 396 653 430 677
rect 396 609 430 615
rect 396 581 430 609
rect 396 541 430 543
rect 396 509 430 541
rect 396 439 430 471
rect 396 437 430 439
rect 396 371 430 399
rect 396 365 430 371
rect 396 303 430 327
rect 396 293 430 303
rect 396 235 430 255
rect 396 221 430 235
rect 488 745 522 759
rect 488 725 522 745
rect 488 677 522 687
rect 488 653 522 677
rect 488 609 522 615
rect 488 581 522 609
rect 488 541 522 543
rect 488 509 522 541
rect 488 439 522 471
rect 488 437 522 439
rect 488 371 522 399
rect 488 365 522 371
rect 488 303 522 327
rect 488 293 522 303
rect 488 235 522 255
rect 488 221 522 235
rect 580 745 614 759
rect 580 725 614 745
rect 580 677 614 687
rect 580 653 614 677
rect 580 609 614 615
rect 580 581 614 609
rect 580 541 614 543
rect 580 509 614 541
rect 580 439 614 471
rect 580 437 614 439
rect 580 371 614 399
rect 580 365 614 371
rect 580 303 614 327
rect 580 293 614 303
rect 580 235 614 255
rect 580 221 614 235
rect 732 745 734 759
rect 734 745 766 759
rect 732 725 766 745
rect 732 677 734 687
rect 734 677 766 687
rect 732 653 766 677
rect 732 609 734 615
rect 734 609 766 615
rect 732 581 766 609
rect 732 541 734 543
rect 734 541 766 543
rect 732 509 766 541
rect 732 439 766 471
rect 732 437 734 439
rect 734 437 766 439
rect 732 371 766 399
rect 732 365 734 371
rect 734 365 766 371
rect 732 303 766 327
rect 732 293 734 303
rect 734 293 766 303
rect 732 235 766 255
rect 732 221 734 235
rect 734 221 766 235
rect 252 123 574 125
rect 252 21 260 123
rect 260 21 566 123
rect 566 21 574 123
rect 252 19 574 21
<< metal1 >>
rect 236 961 590 980
rect 236 855 252 961
rect 574 855 590 961
rect 236 843 590 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 203 759 255 771
rect 203 725 212 759
rect 246 725 255 759
rect 203 687 255 725
rect 203 653 212 687
rect 246 653 255 687
rect 203 615 255 653
rect 203 581 212 615
rect 246 581 255 615
rect 203 543 255 581
rect 203 509 212 543
rect 246 509 255 543
rect 203 471 255 509
rect 203 459 212 471
rect 246 459 255 471
rect 203 399 255 407
rect 203 395 212 399
rect 246 395 255 399
rect 203 331 255 343
rect 203 267 255 279
rect 203 209 255 215
rect 295 765 347 771
rect 295 701 347 713
rect 295 637 347 649
rect 295 581 304 585
rect 338 581 347 585
rect 295 573 347 581
rect 295 509 304 521
rect 338 509 347 521
rect 295 471 347 509
rect 295 437 304 471
rect 338 437 347 471
rect 295 399 347 437
rect 295 365 304 399
rect 338 365 347 399
rect 295 327 347 365
rect 295 293 304 327
rect 338 293 347 327
rect 295 255 347 293
rect 295 221 304 255
rect 338 221 347 255
rect 295 209 347 221
rect 387 759 439 771
rect 387 725 396 759
rect 430 725 439 759
rect 387 687 439 725
rect 387 653 396 687
rect 430 653 439 687
rect 387 615 439 653
rect 387 581 396 615
rect 430 581 439 615
rect 387 543 439 581
rect 387 509 396 543
rect 430 509 439 543
rect 387 471 439 509
rect 387 459 396 471
rect 430 459 439 471
rect 387 399 439 407
rect 387 395 396 399
rect 430 395 439 399
rect 387 331 439 343
rect 387 267 439 279
rect 387 209 439 215
rect 479 765 531 771
rect 479 701 531 713
rect 479 637 531 649
rect 479 581 488 585
rect 522 581 531 585
rect 479 573 531 581
rect 479 509 488 521
rect 522 509 531 521
rect 479 471 531 509
rect 479 437 488 471
rect 522 437 531 471
rect 479 399 531 437
rect 479 365 488 399
rect 522 365 531 399
rect 479 327 531 365
rect 479 293 488 327
rect 522 293 531 327
rect 479 255 531 293
rect 479 221 488 255
rect 522 221 531 255
rect 479 209 531 221
rect 571 759 623 771
rect 571 725 580 759
rect 614 725 623 759
rect 571 687 623 725
rect 571 653 580 687
rect 614 653 623 687
rect 571 615 623 653
rect 571 581 580 615
rect 614 581 623 615
rect 571 543 623 581
rect 571 509 580 543
rect 614 509 623 543
rect 571 471 623 509
rect 571 459 580 471
rect 614 459 623 471
rect 571 399 623 407
rect 571 395 580 399
rect 614 395 623 399
rect 571 331 623 343
rect 571 267 623 279
rect 571 209 623 215
rect 726 759 785 771
rect 726 725 732 759
rect 766 725 785 759
rect 726 687 785 725
rect 726 653 732 687
rect 766 653 785 687
rect 726 615 785 653
rect 726 581 732 615
rect 766 581 785 615
rect 726 543 785 581
rect 726 509 732 543
rect 766 509 785 543
rect 726 471 785 509
rect 726 437 732 471
rect 766 437 785 471
rect 726 399 785 437
rect 726 365 732 399
rect 766 365 785 399
rect 726 327 785 365
rect 726 293 732 327
rect 766 293 785 327
rect 726 255 785 293
rect 726 221 732 255
rect 766 221 785 255
rect 726 209 785 221
rect 236 125 590 137
rect 236 19 252 125
rect 574 19 590 125
rect 236 0 590 19
<< via1 >>
rect 203 437 212 459
rect 212 437 246 459
rect 246 437 255 459
rect 203 407 255 437
rect 203 365 212 395
rect 212 365 246 395
rect 246 365 255 395
rect 203 343 255 365
rect 203 327 255 331
rect 203 293 212 327
rect 212 293 246 327
rect 246 293 255 327
rect 203 279 255 293
rect 203 255 255 267
rect 203 221 212 255
rect 212 221 246 255
rect 246 221 255 255
rect 203 215 255 221
rect 295 759 347 765
rect 295 725 304 759
rect 304 725 338 759
rect 338 725 347 759
rect 295 713 347 725
rect 295 687 347 701
rect 295 653 304 687
rect 304 653 338 687
rect 338 653 347 687
rect 295 649 347 653
rect 295 615 347 637
rect 295 585 304 615
rect 304 585 338 615
rect 338 585 347 615
rect 295 543 347 573
rect 295 521 304 543
rect 304 521 338 543
rect 338 521 347 543
rect 387 437 396 459
rect 396 437 430 459
rect 430 437 439 459
rect 387 407 439 437
rect 387 365 396 395
rect 396 365 430 395
rect 430 365 439 395
rect 387 343 439 365
rect 387 327 439 331
rect 387 293 396 327
rect 396 293 430 327
rect 430 293 439 327
rect 387 279 439 293
rect 387 255 439 267
rect 387 221 396 255
rect 396 221 430 255
rect 430 221 439 255
rect 387 215 439 221
rect 479 759 531 765
rect 479 725 488 759
rect 488 725 522 759
rect 522 725 531 759
rect 479 713 531 725
rect 479 687 531 701
rect 479 653 488 687
rect 488 653 522 687
rect 522 653 531 687
rect 479 649 531 653
rect 479 615 531 637
rect 479 585 488 615
rect 488 585 522 615
rect 522 585 531 615
rect 479 543 531 573
rect 479 521 488 543
rect 488 521 522 543
rect 522 521 531 543
rect 571 437 580 459
rect 580 437 614 459
rect 614 437 623 459
rect 571 407 623 437
rect 571 365 580 395
rect 580 365 614 395
rect 614 365 623 395
rect 571 343 623 365
rect 571 327 623 331
rect 571 293 580 327
rect 580 293 614 327
rect 614 293 623 327
rect 571 279 623 293
rect 571 255 623 267
rect 571 221 580 255
rect 580 221 614 255
rect 614 221 623 255
rect 571 215 623 221
<< metal2 >>
rect 14 765 812 771
rect 14 713 295 765
rect 347 713 479 765
rect 531 713 812 765
rect 14 701 812 713
rect 14 649 295 701
rect 347 649 479 701
rect 531 649 812 701
rect 14 637 812 649
rect 14 585 295 637
rect 347 585 479 637
rect 531 585 812 637
rect 14 573 812 585
rect 14 521 295 573
rect 347 521 479 573
rect 531 521 812 573
rect 14 515 812 521
rect 14 459 812 465
rect 14 407 203 459
rect 255 407 387 459
rect 439 407 571 459
rect 623 407 812 459
rect 14 395 812 407
rect 14 343 203 395
rect 255 343 387 395
rect 439 343 571 395
rect 623 343 812 395
rect 14 331 812 343
rect 14 279 203 331
rect 255 279 387 331
rect 439 279 571 331
rect 623 279 812 331
rect 14 267 812 279
rect 14 215 203 267
rect 255 215 387 267
rect 439 215 571 267
rect 623 215 812 267
rect 14 209 812 215
<< labels >>
flabel metal1 s 301 42 535 92 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 301 878 535 928 0 FreeSans 200 0 0 0 GATE
port 2 nsew
flabel metal1 s 41 466 100 496 0 FreeSans 200 90 0 0 BULK
port 4 nsew
flabel metal1 s 726 469 785 499 0 FreeSans 200 90 0 0 BULK
port 4 nsew
flabel comment s 637 488 637 488 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 184 487 184 487 0 FreeSans 180 90 0 0 dummy_poly
flabel comment s 241 490 241 490 0 FreeSans 300 0 0 0 S
flabel comment s 327 490 327 490 0 FreeSans 300 0 0 0 S
flabel comment s 413 490 413 490 0 FreeSans 300 0 0 0 S
flabel comment s 499 490 499 490 0 FreeSans 300 0 0 0 S
flabel comment s 241 490 241 490 0 FreeSans 300 0 0 0 S
flabel comment s 327 490 327 490 0 FreeSans 300 0 0 0 D
flabel comment s 413 490 413 490 0 FreeSans 300 0 0 0 S
flabel comment s 499 490 499 490 0 FreeSans 300 0 0 0 D
flabel comment s 585 490 585 490 0 FreeSans 300 0 0 0 S
flabel metal2 s 14 280 35 408 7 FreeSans 300 180 0 0 SOURCE
port 3 nsew
flabel metal2 s 14 589 35 717 7 FreeSans 300 180 0 0 DRAIN
port 1 nsew
<< properties >>
string GDS_END 9697378
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9676500
string device primitive
<< end >>
