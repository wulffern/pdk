magic
tech sky130A
magscale 1 2
timestamp 1665766018
<< pwell >>
rect 523 817 544 866
<< obsli1 >>
rect 16 1116 1150 1150
rect 16 50 50 1116
rect 1116 50 1150 1116
rect 16 16 1150 50
<< obsm1 >>
rect 0 66 66 1164
rect 94 1102 1164 1164
rect 94 94 122 1102
rect 150 66 178 1074
rect 206 94 234 1102
rect 262 66 290 1074
rect 318 94 346 1102
rect 374 66 402 1074
rect 430 94 458 1102
rect 486 66 514 1074
rect 542 94 570 1102
rect 598 66 626 1074
rect 654 94 682 1102
rect 710 66 738 1074
rect 766 94 794 1102
rect 822 66 850 1074
rect 878 94 906 1102
rect 934 66 962 1074
rect 990 94 1018 1102
rect 1046 66 1074 1074
rect 1102 94 1164 1102
rect 0 0 1164 66
<< obsm2 >>
rect 66 1102 1164 1164
rect 0 1046 1074 1074
rect 0 962 66 1046
rect 1102 1018 1164 1102
rect 94 990 1164 1018
rect 0 934 1074 962
rect 0 850 66 934
rect 1102 906 1164 990
rect 94 878 1164 906
rect 0 822 1074 850
rect 0 738 66 822
rect 1102 794 1164 878
rect 94 766 1164 794
rect 0 710 1074 738
rect 0 626 66 710
rect 1102 682 1164 766
rect 94 654 1164 682
rect 0 598 1074 626
rect 0 514 66 598
rect 1102 570 1164 654
rect 94 542 1164 570
rect 0 486 1074 514
rect 0 402 66 486
rect 1102 458 1164 542
rect 94 430 1164 458
rect 0 374 1074 402
rect 0 290 66 374
rect 1102 346 1164 430
rect 94 318 1164 346
rect 0 262 1074 290
rect 0 178 66 262
rect 1102 234 1164 318
rect 94 206 1164 234
rect 0 150 1074 178
rect 0 66 66 150
rect 1102 122 1164 206
rect 94 94 1164 122
rect 1102 66 1164 94
rect 0 0 1074 66
<< obsm3 >>
rect 66 1086 1180 1180
rect 0 66 66 1026
rect 126 126 186 1086
rect 246 66 306 1026
rect 366 126 426 1086
rect 486 66 546 1026
rect 606 126 666 1086
rect 726 66 786 1026
rect 846 126 906 1086
rect 966 66 1026 1026
rect 1086 66 1180 1086
rect 0 0 1026 66
<< metal4 >>
rect 0 1026 66 1180
rect 126 1086 1180 1180
rect 0 966 1026 1026
rect 0 786 66 966
rect 1086 906 1180 1086
rect 126 846 1180 906
rect 0 726 1026 786
rect 0 546 66 726
rect 1086 666 1180 846
rect 126 606 1180 666
rect 0 486 1026 546
rect 0 306 66 486
rect 1086 426 1180 606
rect 126 366 1180 426
rect 0 246 1026 306
rect 0 66 66 246
rect 1086 186 1180 366
rect 126 126 1180 186
rect 0 0 1180 66
<< labels >>
rlabel metal4 s 0 1026 66 1180 6 C0
port 1 nsew
rlabel metal4 s 0 966 1026 1026 6 C0
port 1 nsew
rlabel metal4 s 0 786 66 966 6 C0
port 1 nsew
rlabel metal4 s 0 726 1026 786 6 C0
port 1 nsew
rlabel metal4 s 0 546 66 726 6 C0
port 1 nsew
rlabel metal4 s 0 486 1026 546 6 C0
port 1 nsew
rlabel metal4 s 0 306 66 486 6 C0
port 1 nsew
rlabel metal4 s 0 246 1026 306 6 C0
port 1 nsew
rlabel metal4 s 0 66 66 246 6 C0
port 1 nsew
rlabel metal4 s 0 0 1180 66 6 C0
port 1 nsew
rlabel metal4 s 1086 906 1180 1086 6 C1
port 2 nsew
rlabel metal4 s 1086 666 1180 846 6 C1
port 2 nsew
rlabel metal4 s 1086 426 1180 606 6 C1
port 2 nsew
rlabel metal4 s 1086 186 1180 366 6 C1
port 2 nsew
rlabel metal4 s 126 1086 1180 1180 6 C1
port 2 nsew
rlabel metal4 s 126 846 1180 906 6 C1
port 2 nsew
rlabel metal4 s 126 606 1180 666 6 C1
port 2 nsew
rlabel metal4 s 126 366 1180 426 6 C1
port 2 nsew
rlabel metal4 s 126 126 1180 186 6 C1
port 2 nsew
rlabel pwell s 523 817 544 866 6 SUB
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 1180 1180
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 169568
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 155424
string device primitive
<< end >>
