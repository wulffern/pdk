/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/corners/ss/specialized_cells.spice