magic
tech sky130A
magscale 1 2
timestamp 1665766018
<< nwell >>
rect 148 604 1052 1896
<< pmos >>
rect 352 745 382 1755
rect 506 745 536 1755
rect 660 745 690 1755
rect 814 745 844 1755
<< pdiff >>
rect 296 1743 352 1755
rect 296 1709 307 1743
rect 341 1709 352 1743
rect 296 1675 352 1709
rect 296 1641 307 1675
rect 341 1641 352 1675
rect 296 1607 352 1641
rect 296 1573 307 1607
rect 341 1573 352 1607
rect 296 1539 352 1573
rect 296 1505 307 1539
rect 341 1505 352 1539
rect 296 1471 352 1505
rect 296 1437 307 1471
rect 341 1437 352 1471
rect 296 1403 352 1437
rect 296 1369 307 1403
rect 341 1369 352 1403
rect 296 1335 352 1369
rect 296 1301 307 1335
rect 341 1301 352 1335
rect 296 1267 352 1301
rect 296 1233 307 1267
rect 341 1233 352 1267
rect 296 1199 352 1233
rect 296 1165 307 1199
rect 341 1165 352 1199
rect 296 1131 352 1165
rect 296 1097 307 1131
rect 341 1097 352 1131
rect 296 1063 352 1097
rect 296 1029 307 1063
rect 341 1029 352 1063
rect 296 995 352 1029
rect 296 961 307 995
rect 341 961 352 995
rect 296 927 352 961
rect 296 893 307 927
rect 341 893 352 927
rect 296 859 352 893
rect 296 825 307 859
rect 341 825 352 859
rect 296 791 352 825
rect 296 757 307 791
rect 341 757 352 791
rect 296 745 352 757
rect 382 1743 506 1755
rect 382 757 393 1743
rect 495 757 506 1743
rect 382 745 506 757
rect 536 1743 660 1755
rect 536 757 547 1743
rect 649 757 660 1743
rect 536 745 660 757
rect 690 1743 814 1755
rect 690 757 701 1743
rect 803 757 814 1743
rect 690 745 814 757
rect 844 1743 903 1755
rect 844 1709 855 1743
rect 889 1709 903 1743
rect 844 1675 903 1709
rect 844 1641 855 1675
rect 889 1641 903 1675
rect 844 1607 903 1641
rect 844 1573 855 1607
rect 889 1573 903 1607
rect 844 1539 903 1573
rect 844 1505 855 1539
rect 889 1505 903 1539
rect 844 1471 903 1505
rect 844 1437 855 1471
rect 889 1437 903 1471
rect 844 1403 903 1437
rect 844 1369 855 1403
rect 889 1369 903 1403
rect 844 1335 903 1369
rect 844 1301 855 1335
rect 889 1301 903 1335
rect 844 1267 903 1301
rect 844 1233 855 1267
rect 889 1233 903 1267
rect 844 1199 903 1233
rect 844 1165 855 1199
rect 889 1165 903 1199
rect 844 1131 903 1165
rect 844 1097 855 1131
rect 889 1097 903 1131
rect 844 1063 903 1097
rect 844 1029 855 1063
rect 889 1029 903 1063
rect 844 995 903 1029
rect 844 961 855 995
rect 889 961 903 995
rect 844 927 903 961
rect 844 893 855 927
rect 889 893 903 927
rect 844 859 903 893
rect 844 825 855 859
rect 889 825 903 859
rect 844 791 903 825
rect 844 757 855 791
rect 889 757 903 791
rect 844 745 903 757
<< pdiffc >>
rect 307 1709 341 1743
rect 307 1641 341 1675
rect 307 1573 341 1607
rect 307 1505 341 1539
rect 307 1437 341 1471
rect 307 1369 341 1403
rect 307 1301 341 1335
rect 307 1233 341 1267
rect 307 1165 341 1199
rect 307 1097 341 1131
rect 307 1029 341 1063
rect 307 961 341 995
rect 307 893 341 927
rect 307 825 341 859
rect 307 757 341 791
rect 393 757 495 1743
rect 547 757 649 1743
rect 701 757 803 1743
rect 855 1709 889 1743
rect 855 1641 889 1675
rect 855 1573 889 1607
rect 855 1505 889 1539
rect 855 1437 889 1471
rect 855 1369 889 1403
rect 855 1301 889 1335
rect 855 1233 889 1267
rect 855 1165 889 1199
rect 855 1097 889 1131
rect 855 1029 889 1063
rect 855 961 889 995
rect 855 893 889 927
rect 855 825 889 859
rect 855 757 889 791
<< nsubdiff >>
rect 184 1709 242 1755
rect 184 1675 196 1709
rect 230 1675 242 1709
rect 184 1641 242 1675
rect 184 1607 196 1641
rect 230 1607 242 1641
rect 184 1573 242 1607
rect 184 1539 196 1573
rect 230 1539 242 1573
rect 184 1505 242 1539
rect 184 1471 196 1505
rect 230 1471 242 1505
rect 184 1437 242 1471
rect 184 1403 196 1437
rect 230 1403 242 1437
rect 184 1369 242 1403
rect 184 1335 196 1369
rect 230 1335 242 1369
rect 184 1301 242 1335
rect 184 1267 196 1301
rect 230 1267 242 1301
rect 184 1233 242 1267
rect 184 1199 196 1233
rect 230 1199 242 1233
rect 184 1165 242 1199
rect 184 1131 196 1165
rect 230 1131 242 1165
rect 184 1097 242 1131
rect 184 1063 196 1097
rect 230 1063 242 1097
rect 184 1029 242 1063
rect 184 995 196 1029
rect 230 995 242 1029
rect 184 961 242 995
rect 184 927 196 961
rect 230 927 242 961
rect 184 893 242 927
rect 184 859 196 893
rect 230 859 242 893
rect 184 825 242 859
rect 184 791 196 825
rect 230 791 242 825
rect 184 745 242 791
rect 957 1709 1015 1755
rect 957 1675 969 1709
rect 1003 1675 1015 1709
rect 957 1641 1015 1675
rect 957 1607 969 1641
rect 1003 1607 1015 1641
rect 957 1573 1015 1607
rect 957 1539 969 1573
rect 1003 1539 1015 1573
rect 957 1505 1015 1539
rect 957 1471 969 1505
rect 1003 1471 1015 1505
rect 957 1437 1015 1471
rect 957 1403 969 1437
rect 1003 1403 1015 1437
rect 957 1369 1015 1403
rect 957 1335 969 1369
rect 1003 1335 1015 1369
rect 957 1301 1015 1335
rect 957 1267 969 1301
rect 1003 1267 1015 1301
rect 957 1233 1015 1267
rect 957 1199 969 1233
rect 1003 1199 1015 1233
rect 957 1165 1015 1199
rect 957 1131 969 1165
rect 1003 1131 1015 1165
rect 957 1097 1015 1131
rect 957 1063 969 1097
rect 1003 1063 1015 1097
rect 957 1029 1015 1063
rect 957 995 969 1029
rect 1003 995 1015 1029
rect 957 961 1015 995
rect 957 927 969 961
rect 1003 927 1015 961
rect 957 893 1015 927
rect 957 859 969 893
rect 1003 859 1015 893
rect 957 825 1015 859
rect 957 791 969 825
rect 1003 791 1015 825
rect 957 745 1015 791
<< nsubdiffcont >>
rect 196 1675 230 1709
rect 196 1607 230 1641
rect 196 1539 230 1573
rect 196 1471 230 1505
rect 196 1403 230 1437
rect 196 1335 230 1369
rect 196 1267 230 1301
rect 196 1199 230 1233
rect 196 1131 230 1165
rect 196 1063 230 1097
rect 196 995 230 1029
rect 196 927 230 961
rect 196 859 230 893
rect 196 791 230 825
rect 969 1675 1003 1709
rect 969 1607 1003 1641
rect 969 1539 1003 1573
rect 969 1471 1003 1505
rect 969 1403 1003 1437
rect 969 1335 1003 1369
rect 969 1267 1003 1301
rect 969 1199 1003 1233
rect 969 1131 1003 1165
rect 969 1063 1003 1097
rect 969 995 1003 1029
rect 969 927 1003 961
rect 969 859 1003 893
rect 969 791 1003 825
<< poly >>
rect 352 1850 894 1866
rect 352 1816 368 1850
rect 402 1816 436 1850
rect 470 1816 504 1850
rect 538 1816 572 1850
rect 606 1816 640 1850
rect 674 1816 708 1850
rect 742 1816 776 1850
rect 810 1816 844 1850
rect 878 1816 894 1850
rect 352 1800 894 1816
rect 352 1755 382 1800
rect 506 1755 536 1800
rect 660 1755 690 1800
rect 814 1755 844 1800
rect 352 700 382 745
rect 506 700 536 745
rect 660 700 690 745
rect 814 700 844 745
rect 352 684 894 700
rect 352 650 368 684
rect 402 650 436 684
rect 470 650 504 684
rect 538 650 572 684
rect 606 650 640 684
rect 674 650 708 684
rect 742 650 776 684
rect 810 650 844 684
rect 878 650 894 684
rect 352 634 894 650
<< polycont >>
rect 368 1816 402 1850
rect 436 1816 470 1850
rect 504 1816 538 1850
rect 572 1816 606 1850
rect 640 1816 674 1850
rect 708 1816 742 1850
rect 776 1816 810 1850
rect 844 1816 878 1850
rect 368 650 402 684
rect 436 650 470 684
rect 504 650 538 684
rect 572 650 606 684
rect 640 650 674 684
rect 708 650 742 684
rect 776 650 810 684
rect 844 650 878 684
<< locali >>
rect 402 1816 424 1850
rect 470 1816 496 1850
rect 538 1816 568 1850
rect 606 1816 640 1850
rect 674 1816 708 1850
rect 746 1816 776 1850
rect 818 1816 844 1850
rect 890 1816 894 1850
rect 307 1743 341 1759
rect 196 1663 230 1675
rect 196 1591 230 1607
rect 196 1519 230 1539
rect 196 1447 230 1471
rect 196 1375 230 1403
rect 196 1303 230 1335
rect 196 1233 230 1267
rect 196 1165 230 1197
rect 196 1097 230 1125
rect 196 1029 230 1053
rect 196 961 230 981
rect 196 893 230 909
rect 196 825 230 837
rect 307 1675 341 1701
rect 307 1607 341 1629
rect 307 1539 341 1557
rect 307 1471 341 1485
rect 307 1403 341 1413
rect 307 1335 341 1341
rect 307 1267 341 1269
rect 307 1231 341 1233
rect 307 1159 341 1165
rect 307 1087 341 1097
rect 307 1015 341 1029
rect 307 943 341 961
rect 307 871 341 893
rect 307 799 341 825
rect 307 741 341 757
rect 391 1743 497 1759
rect 391 1735 393 1743
rect 495 1735 497 1743
rect 391 757 393 765
rect 495 757 497 765
rect 391 741 497 757
rect 545 1743 651 1759
rect 545 1735 547 1743
rect 649 1735 651 1743
rect 545 757 547 765
rect 649 757 651 765
rect 545 741 651 757
rect 699 1743 805 1759
rect 699 1735 701 1743
rect 803 1735 805 1743
rect 699 757 701 765
rect 803 757 805 765
rect 699 741 805 757
rect 855 1743 889 1759
rect 855 1675 889 1701
rect 855 1607 889 1629
rect 855 1539 889 1557
rect 855 1471 889 1485
rect 855 1403 889 1413
rect 855 1335 889 1341
rect 855 1267 889 1269
rect 855 1231 889 1233
rect 855 1159 889 1165
rect 855 1087 889 1097
rect 855 1015 889 1029
rect 855 943 889 961
rect 855 871 889 893
rect 855 799 889 825
rect 969 1663 1003 1675
rect 969 1591 1003 1607
rect 969 1519 1003 1539
rect 969 1447 1003 1471
rect 969 1375 1003 1403
rect 969 1303 1003 1335
rect 969 1233 1003 1267
rect 969 1165 1003 1197
rect 969 1097 1003 1125
rect 969 1029 1003 1053
rect 969 961 1003 981
rect 969 893 1003 909
rect 969 825 1003 837
rect 855 741 889 757
rect 402 650 424 684
rect 470 650 496 684
rect 538 650 568 684
rect 606 650 640 684
rect 674 650 708 684
rect 746 650 776 684
rect 818 650 844 684
rect 890 650 894 684
<< viali >>
rect 352 1816 368 1850
rect 368 1816 386 1850
rect 424 1816 436 1850
rect 436 1816 458 1850
rect 496 1816 504 1850
rect 504 1816 530 1850
rect 568 1816 572 1850
rect 572 1816 602 1850
rect 640 1816 674 1850
rect 712 1816 742 1850
rect 742 1816 746 1850
rect 784 1816 810 1850
rect 810 1816 818 1850
rect 856 1816 878 1850
rect 878 1816 890 1850
rect 196 1709 230 1735
rect 196 1701 230 1709
rect 196 1641 230 1663
rect 196 1629 230 1641
rect 196 1573 230 1591
rect 196 1557 230 1573
rect 196 1505 230 1519
rect 196 1485 230 1505
rect 196 1437 230 1447
rect 196 1413 230 1437
rect 196 1369 230 1375
rect 196 1341 230 1369
rect 196 1301 230 1303
rect 196 1269 230 1301
rect 196 1199 230 1231
rect 196 1197 230 1199
rect 196 1131 230 1159
rect 196 1125 230 1131
rect 196 1063 230 1087
rect 196 1053 230 1063
rect 196 995 230 1015
rect 196 981 230 995
rect 196 927 230 943
rect 196 909 230 927
rect 196 859 230 871
rect 196 837 230 859
rect 196 791 230 799
rect 196 765 230 791
rect 307 1709 341 1735
rect 307 1701 341 1709
rect 307 1641 341 1663
rect 307 1629 341 1641
rect 307 1573 341 1591
rect 307 1557 341 1573
rect 307 1505 341 1519
rect 307 1485 341 1505
rect 307 1437 341 1447
rect 307 1413 341 1437
rect 307 1369 341 1375
rect 307 1341 341 1369
rect 307 1301 341 1303
rect 307 1269 341 1301
rect 307 1199 341 1231
rect 307 1197 341 1199
rect 307 1131 341 1159
rect 307 1125 341 1131
rect 307 1063 341 1087
rect 307 1053 341 1063
rect 307 995 341 1015
rect 307 981 341 995
rect 307 927 341 943
rect 307 909 341 927
rect 307 859 341 871
rect 307 837 341 859
rect 307 791 341 799
rect 307 765 341 791
rect 391 765 393 1735
rect 393 765 495 1735
rect 495 765 497 1735
rect 545 765 547 1735
rect 547 765 649 1735
rect 649 765 651 1735
rect 699 765 701 1735
rect 701 765 803 1735
rect 803 765 805 1735
rect 855 1709 889 1735
rect 855 1701 889 1709
rect 855 1641 889 1663
rect 855 1629 889 1641
rect 855 1573 889 1591
rect 855 1557 889 1573
rect 855 1505 889 1519
rect 855 1485 889 1505
rect 855 1437 889 1447
rect 855 1413 889 1437
rect 855 1369 889 1375
rect 855 1341 889 1369
rect 855 1301 889 1303
rect 855 1269 889 1301
rect 855 1199 889 1231
rect 855 1197 889 1199
rect 855 1131 889 1159
rect 855 1125 889 1131
rect 855 1063 889 1087
rect 855 1053 889 1063
rect 855 995 889 1015
rect 855 981 889 995
rect 855 927 889 943
rect 855 909 889 927
rect 855 859 889 871
rect 855 837 889 859
rect 855 791 889 799
rect 855 765 889 791
rect 969 1709 1003 1735
rect 969 1701 1003 1709
rect 969 1641 1003 1663
rect 969 1629 1003 1641
rect 969 1573 1003 1591
rect 969 1557 1003 1573
rect 969 1505 1003 1519
rect 969 1485 1003 1505
rect 969 1437 1003 1447
rect 969 1413 1003 1437
rect 969 1369 1003 1375
rect 969 1341 1003 1369
rect 969 1301 1003 1303
rect 969 1269 1003 1301
rect 969 1199 1003 1231
rect 969 1197 1003 1199
rect 969 1131 1003 1159
rect 969 1125 1003 1131
rect 969 1063 1003 1087
rect 969 1053 1003 1063
rect 969 995 1003 1015
rect 969 981 1003 995
rect 969 927 1003 943
rect 969 909 1003 927
rect 969 859 1003 871
rect 969 837 1003 859
rect 969 791 1003 799
rect 969 765 1003 791
rect 352 650 368 684
rect 368 650 386 684
rect 424 650 436 684
rect 436 650 458 684
rect 496 650 504 684
rect 504 650 530 684
rect 568 650 572 684
rect 572 650 602 684
rect 640 650 674 684
rect 712 650 742 684
rect 742 650 746 684
rect 784 650 810 684
rect 810 650 818 684
rect 856 650 878 684
rect 878 650 890 684
<< metal1 >>
rect 340 1850 902 1862
rect 340 1816 352 1850
rect 386 1816 424 1850
rect 458 1816 496 1850
rect 530 1816 568 1850
rect 602 1816 640 1850
rect 674 1816 712 1850
rect 746 1816 784 1850
rect 818 1816 856 1850
rect 890 1816 902 1850
rect 340 1804 902 1816
rect 298 1770 350 1776
rect 184 1735 242 1747
rect 184 1701 196 1735
rect 230 1701 242 1735
rect 184 1663 242 1701
rect 184 1629 196 1663
rect 230 1629 242 1663
rect 184 1591 242 1629
rect 184 1557 196 1591
rect 230 1557 242 1591
rect 184 1519 242 1557
rect 184 1485 196 1519
rect 230 1485 242 1519
rect 184 1447 242 1485
rect 184 1413 196 1447
rect 230 1413 242 1447
rect 184 1375 242 1413
rect 184 1341 196 1375
rect 230 1341 242 1375
rect 184 1303 242 1341
rect 184 1269 196 1303
rect 230 1269 242 1303
rect 184 1231 242 1269
rect 184 1197 196 1231
rect 230 1197 242 1231
rect 184 1159 242 1197
rect 184 1125 196 1159
rect 230 1125 242 1159
rect 184 1087 242 1125
rect 184 1053 196 1087
rect 230 1053 242 1087
rect 184 1015 242 1053
rect 184 981 196 1015
rect 230 981 242 1015
rect 184 943 242 981
rect 184 909 196 943
rect 230 909 242 943
rect 184 871 242 909
rect 184 837 196 871
rect 230 837 242 871
rect 184 799 242 837
rect 184 765 196 799
rect 230 765 242 799
rect 184 753 242 765
rect 540 1770 656 1776
rect 350 1718 353 1747
rect 298 1706 307 1718
rect 341 1706 353 1718
rect 350 1654 353 1706
rect 298 1642 307 1654
rect 341 1642 353 1654
rect 350 1590 353 1642
rect 298 1578 307 1590
rect 341 1578 353 1590
rect 350 1526 353 1578
rect 298 1519 353 1526
rect 298 1514 307 1519
rect 341 1514 353 1519
rect 350 1462 353 1514
rect 298 1447 353 1462
rect 298 1413 307 1447
rect 341 1413 353 1447
rect 298 1375 353 1413
rect 298 1341 307 1375
rect 341 1341 353 1375
rect 298 1303 353 1341
rect 298 1269 307 1303
rect 341 1269 353 1303
rect 298 1231 353 1269
rect 298 1197 307 1231
rect 341 1197 353 1231
rect 298 1159 353 1197
rect 298 1125 307 1159
rect 341 1125 353 1159
rect 298 1087 353 1125
rect 298 1053 307 1087
rect 341 1053 353 1087
rect 298 1038 353 1053
rect 350 986 353 1038
rect 298 981 307 986
rect 341 981 353 986
rect 298 974 353 981
rect 350 922 353 974
rect 298 910 307 922
rect 341 910 353 922
rect 350 858 353 910
rect 298 846 307 858
rect 341 846 353 858
rect 350 794 353 846
rect 298 782 307 794
rect 341 782 353 794
rect 350 753 353 782
rect 381 1735 507 1747
rect 381 1564 391 1735
rect 497 1564 507 1735
rect 381 936 386 1564
rect 502 936 507 1564
rect 381 765 391 936
rect 497 765 507 936
rect 381 753 507 765
rect 535 1462 540 1747
rect 846 1770 898 1776
rect 656 1462 661 1747
rect 535 1038 545 1462
rect 651 1038 661 1462
rect 535 753 540 1038
rect 298 724 350 730
rect 656 753 661 1038
rect 689 1735 815 1747
rect 689 1564 699 1735
rect 805 1564 815 1735
rect 689 936 694 1564
rect 810 936 815 1564
rect 689 765 699 936
rect 805 765 815 936
rect 689 753 815 765
rect 843 1718 846 1747
rect 898 1718 901 1747
rect 843 1706 855 1718
rect 889 1706 901 1718
rect 843 1654 846 1706
rect 898 1654 901 1706
rect 843 1642 855 1654
rect 889 1642 901 1654
rect 843 1590 846 1642
rect 898 1590 901 1642
rect 843 1578 855 1590
rect 889 1578 901 1590
rect 843 1526 846 1578
rect 898 1526 901 1578
rect 843 1519 901 1526
rect 843 1514 855 1519
rect 889 1514 901 1519
rect 843 1462 846 1514
rect 898 1462 901 1514
rect 843 1447 901 1462
rect 843 1413 855 1447
rect 889 1413 901 1447
rect 843 1375 901 1413
rect 843 1341 855 1375
rect 889 1341 901 1375
rect 843 1303 901 1341
rect 843 1269 855 1303
rect 889 1269 901 1303
rect 843 1231 901 1269
rect 843 1197 855 1231
rect 889 1197 901 1231
rect 843 1159 901 1197
rect 843 1125 855 1159
rect 889 1125 901 1159
rect 843 1087 901 1125
rect 843 1053 855 1087
rect 889 1053 901 1087
rect 843 1038 901 1053
rect 843 986 846 1038
rect 898 986 901 1038
rect 843 981 855 986
rect 889 981 901 986
rect 843 974 901 981
rect 843 922 846 974
rect 898 922 901 974
rect 843 910 855 922
rect 889 910 901 922
rect 843 858 846 910
rect 898 858 901 910
rect 843 846 855 858
rect 889 846 901 858
rect 843 794 846 846
rect 898 794 901 846
rect 843 782 855 794
rect 889 782 901 794
rect 843 753 846 782
rect 540 724 656 730
rect 898 753 901 782
rect 957 1735 1015 1747
rect 957 1701 969 1735
rect 1003 1701 1015 1735
rect 957 1663 1015 1701
rect 957 1629 969 1663
rect 1003 1629 1015 1663
rect 957 1591 1015 1629
rect 957 1557 969 1591
rect 1003 1557 1015 1591
rect 957 1519 1015 1557
rect 957 1485 969 1519
rect 1003 1485 1015 1519
rect 957 1447 1015 1485
rect 957 1413 969 1447
rect 1003 1413 1015 1447
rect 957 1375 1015 1413
rect 957 1341 969 1375
rect 1003 1341 1015 1375
rect 957 1303 1015 1341
rect 957 1269 969 1303
rect 1003 1269 1015 1303
rect 957 1231 1015 1269
rect 957 1197 969 1231
rect 1003 1197 1015 1231
rect 957 1159 1015 1197
rect 957 1125 969 1159
rect 1003 1125 1015 1159
rect 957 1087 1015 1125
rect 957 1053 969 1087
rect 1003 1053 1015 1087
rect 957 1015 1015 1053
rect 957 981 969 1015
rect 1003 981 1015 1015
rect 957 943 1015 981
rect 957 909 969 943
rect 1003 909 1015 943
rect 957 871 1015 909
rect 957 837 969 871
rect 1003 837 1015 871
rect 957 799 1015 837
rect 957 765 969 799
rect 1003 765 1015 799
rect 957 753 1015 765
rect 846 724 898 730
rect 340 684 902 696
rect 340 650 352 684
rect 386 650 424 684
rect 458 650 496 684
rect 530 650 568 684
rect 602 650 640 684
rect 674 650 712 684
rect 746 650 784 684
rect 818 650 856 684
rect 890 650 902 684
rect 340 638 902 650
<< via1 >>
rect 298 1735 350 1770
rect 298 1718 307 1735
rect 307 1718 341 1735
rect 341 1718 350 1735
rect 298 1701 307 1706
rect 307 1701 341 1706
rect 341 1701 350 1706
rect 298 1663 350 1701
rect 298 1654 307 1663
rect 307 1654 341 1663
rect 341 1654 350 1663
rect 298 1629 307 1642
rect 307 1629 341 1642
rect 341 1629 350 1642
rect 298 1591 350 1629
rect 298 1590 307 1591
rect 307 1590 341 1591
rect 341 1590 350 1591
rect 298 1557 307 1578
rect 307 1557 341 1578
rect 341 1557 350 1578
rect 298 1526 350 1557
rect 298 1485 307 1514
rect 307 1485 341 1514
rect 341 1485 350 1514
rect 298 1462 350 1485
rect 298 1015 350 1038
rect 298 986 307 1015
rect 307 986 341 1015
rect 341 986 350 1015
rect 298 943 350 974
rect 298 922 307 943
rect 307 922 341 943
rect 341 922 350 943
rect 298 909 307 910
rect 307 909 341 910
rect 341 909 350 910
rect 298 871 350 909
rect 298 858 307 871
rect 307 858 341 871
rect 341 858 350 871
rect 298 837 307 846
rect 307 837 341 846
rect 341 837 350 846
rect 298 799 350 837
rect 298 794 307 799
rect 307 794 341 799
rect 341 794 350 799
rect 298 765 307 782
rect 307 765 341 782
rect 341 765 350 782
rect 298 730 350 765
rect 386 936 391 1564
rect 391 936 497 1564
rect 497 936 502 1564
rect 540 1735 656 1770
rect 540 1462 545 1735
rect 545 1462 651 1735
rect 651 1462 656 1735
rect 540 765 545 1038
rect 545 765 651 1038
rect 651 765 656 1038
rect 540 730 656 765
rect 694 936 699 1564
rect 699 936 805 1564
rect 805 936 810 1564
rect 846 1735 898 1770
rect 846 1718 855 1735
rect 855 1718 889 1735
rect 889 1718 898 1735
rect 846 1701 855 1706
rect 855 1701 889 1706
rect 889 1701 898 1706
rect 846 1663 898 1701
rect 846 1654 855 1663
rect 855 1654 889 1663
rect 889 1654 898 1663
rect 846 1629 855 1642
rect 855 1629 889 1642
rect 889 1629 898 1642
rect 846 1591 898 1629
rect 846 1590 855 1591
rect 855 1590 889 1591
rect 889 1590 898 1591
rect 846 1557 855 1578
rect 855 1557 889 1578
rect 889 1557 898 1578
rect 846 1526 898 1557
rect 846 1485 855 1514
rect 855 1485 889 1514
rect 889 1485 898 1514
rect 846 1462 898 1485
rect 846 1015 898 1038
rect 846 986 855 1015
rect 855 986 889 1015
rect 889 986 898 1015
rect 846 943 898 974
rect 846 922 855 943
rect 855 922 889 943
rect 889 922 898 943
rect 846 909 855 910
rect 855 909 889 910
rect 889 909 898 910
rect 846 871 898 909
rect 846 858 855 871
rect 855 858 889 871
rect 889 858 898 871
rect 846 837 855 846
rect 855 837 889 846
rect 889 837 898 846
rect 846 799 898 837
rect 846 794 855 799
rect 855 794 889 799
rect 889 794 898 799
rect 846 765 855 782
rect 855 765 889 782
rect 889 765 898 782
rect 846 730 898 765
<< metal2 >>
rect 158 2378 1042 2428
rect 158 2122 470 2378
rect 726 2122 1042 2378
rect 158 1770 1042 2122
rect 158 1718 298 1770
rect 350 1718 540 1770
rect 158 1706 540 1718
rect 158 1654 298 1706
rect 350 1654 540 1706
rect 158 1642 540 1654
rect 158 1590 298 1642
rect 350 1626 540 1642
rect 158 1578 350 1590
rect 158 1526 298 1578
rect 158 1514 350 1526
rect 158 1462 298 1514
rect 158 1456 350 1462
rect 386 1564 502 1570
rect 158 1044 214 1456
rect 656 1718 846 1770
rect 898 1718 1042 1770
rect 656 1706 1042 1718
rect 656 1654 846 1706
rect 898 1654 1042 1706
rect 656 1642 1042 1654
rect 656 1626 846 1642
rect 898 1590 1042 1642
rect 846 1578 1042 1590
rect 540 1456 656 1462
rect 694 1564 810 1570
rect 502 1378 694 1428
rect 898 1526 1042 1578
rect 846 1514 1042 1526
rect 898 1462 1042 1514
rect 846 1456 1042 1462
rect 158 1038 350 1044
rect 158 986 298 1038
rect 158 974 350 986
rect 158 922 298 974
rect 502 1072 694 1122
rect 386 930 502 936
rect 540 1038 656 1044
rect 158 910 350 922
rect 158 858 298 910
rect 350 858 540 874
rect 158 846 540 858
rect 158 794 298 846
rect 350 794 540 846
rect 158 782 540 794
rect 158 730 298 782
rect 350 730 540 782
rect 986 1044 1042 1456
rect 694 930 810 936
rect 846 1038 1042 1044
rect 898 986 1042 1038
rect 846 974 1042 986
rect 898 922 1042 974
rect 846 910 1042 922
rect 656 858 846 874
rect 898 858 1042 910
rect 656 846 1042 858
rect 656 794 846 846
rect 898 794 1042 846
rect 656 782 1042 794
rect 656 730 846 782
rect 898 730 1042 782
rect 158 378 1042 730
rect 158 122 470 378
rect 726 122 1042 378
rect 158 72 1042 122
<< via2 >>
rect 470 2122 726 2378
rect 470 1122 502 1378
rect 502 1122 694 1378
rect 694 1122 726 1378
rect 470 122 726 378
<< metal3 >>
rect 0 2378 1200 2500
rect 0 2122 470 2378
rect 726 2122 1200 2378
rect 0 2000 1200 2122
rect 0 1378 1200 1500
rect 0 1122 470 1378
rect 726 1122 1200 1378
rect 0 1000 1200 1122
rect 0 378 1200 500
rect 0 122 470 378
rect 726 122 1200 378
rect 0 0 1200 122
<< labels >>
flabel comment s 436 1285 436 1285 0 FreeSans 300 0 0 0 D
flabel comment s 895 1285 895 1285 0 FreeSans 300 0 0 0 S
flabel comment s 590 1285 590 1285 0 FreeSans 300 0 0 0 S
flabel comment s 316 1285 316 1285 0 FreeSans 300 180 0 0 S
flabel comment s 744 1285 744 1285 0 FreeSans 300 0 0 0 D
flabel metal2 s 430 963 459 1036 0 FreeSans 200 0 0 0 DRAIN
port 1 nsew
flabel metal2 s 203 1786 232 1859 0 FreeSans 200 0 0 0 SOURCE
port 2 nsew
flabel metal1 s 559 653 632 682 0 FreeSans 200 90 0 0 GATE
port 3 nsew
flabel metal1 s 203 1231 232 1304 0 FreeSans 200 0 0 0 BULK
port 4 nsew
<< properties >>
string GDS_END 9881838
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9849760
<< end >>
