/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/corners/ss/rf.spice