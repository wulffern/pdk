/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__esd_rf_nfet_20v0_iec_21vW60p00.spice