/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_see_e/begin_of_life/typical.spice