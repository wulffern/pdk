/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__cap_vpp_33p6x23p1_pol1m1m2m3m4m5_noshield.spice