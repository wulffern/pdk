/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/r+c/res_low__cap_low__lin.spice