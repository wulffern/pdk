/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_see_p/begin_of_life.pm3.spice