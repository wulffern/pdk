magic
tech sky130B
magscale 1 2
timestamp 1665766018
<< pwell >>
rect -13 -26 73 4246
rect 255 566 276 615
rect 467 -26 553 4246
<< locali >>
rect 13 0 47 4220
rect 493 0 527 4220
<< metal1 >>
rect 14 4213 526 4220
rect 14 4161 44 4213
rect 96 4161 284 4213
rect 336 4161 364 4213
rect 416 4161 444 4213
rect 496 4161 526 4213
rect 14 4154 526 4161
rect 14 126 46 4154
rect 74 66 106 4094
rect 134 126 166 4154
rect 194 66 226 4094
rect 254 126 286 4154
rect 314 66 346 4094
rect 374 126 406 4154
rect 434 66 466 4094
rect 494 126 526 4154
rect 60 59 480 66
rect 60 7 84 59
rect 136 7 164 59
rect 216 7 244 59
rect 296 7 324 59
rect 376 7 404 59
rect 456 7 480 59
rect 60 0 480 7
<< via1 >>
rect 44 4161 96 4213
rect 284 4161 336 4213
rect 364 4161 416 4213
rect 444 4161 496 4213
rect 84 7 136 59
rect 164 7 216 59
rect 244 7 296 59
rect 324 7 376 59
rect 404 7 456 59
<< metal2 >>
rect 14 4215 166 4220
rect 14 4159 42 4215
rect 98 4159 166 4215
rect 14 4154 166 4159
rect 14 126 46 4154
rect 74 66 106 4094
rect 134 126 166 4154
rect 194 66 226 4220
rect 254 4215 526 4220
rect 254 4159 282 4215
rect 338 4159 362 4215
rect 418 4159 442 4215
rect 498 4159 526 4215
rect 254 4154 526 4159
rect 254 126 286 4154
rect 314 66 346 4094
rect 374 126 406 4154
rect 434 66 466 4094
rect 494 126 526 4154
rect 60 61 480 66
rect 60 5 82 61
rect 138 5 162 61
rect 218 5 242 61
rect 298 5 322 61
rect 378 5 402 61
rect 458 5 480 61
rect 60 0 480 5
<< via2 >>
rect 42 4213 98 4215
rect 42 4161 44 4213
rect 44 4161 96 4213
rect 96 4161 98 4213
rect 42 4159 98 4161
rect 282 4213 338 4215
rect 282 4161 284 4213
rect 284 4161 336 4213
rect 336 4161 338 4213
rect 282 4159 338 4161
rect 362 4213 418 4215
rect 362 4161 364 4213
rect 364 4161 416 4213
rect 416 4161 418 4213
rect 362 4159 418 4161
rect 442 4213 498 4215
rect 442 4161 444 4213
rect 444 4161 496 4213
rect 496 4161 498 4213
rect 442 4159 498 4161
rect 82 59 138 61
rect 82 7 84 59
rect 84 7 136 59
rect 136 7 138 59
rect 82 5 138 7
rect 162 59 218 61
rect 162 7 164 59
rect 164 7 216 59
rect 216 7 218 59
rect 162 5 218 7
rect 242 59 298 61
rect 242 7 244 59
rect 244 7 296 59
rect 296 7 298 59
rect 242 5 298 7
rect 322 59 378 61
rect 322 7 324 59
rect 324 7 376 59
rect 376 7 378 59
rect 322 5 378 7
rect 402 59 458 61
rect 402 7 404 59
rect 404 7 456 59
rect 456 7 458 59
rect 402 5 458 7
<< metal3 >>
rect 0 4219 540 4220
rect 0 4155 38 4219
rect 102 4155 118 4219
rect 182 4155 198 4219
rect 262 4155 278 4219
rect 342 4155 358 4219
rect 422 4155 438 4219
rect 502 4155 540 4219
rect 0 4154 540 4155
rect 0 126 60 4154
rect 120 66 180 4094
rect 240 126 300 4154
rect 360 66 420 4094
rect 480 126 540 4154
rect 60 65 480 66
rect 60 1 78 65
rect 142 1 158 65
rect 222 1 238 65
rect 302 1 318 65
rect 382 1 398 65
rect 462 1 480 65
rect 60 0 480 1
<< via3 >>
rect 38 4215 102 4219
rect 38 4159 42 4215
rect 42 4159 98 4215
rect 98 4159 102 4215
rect 38 4155 102 4159
rect 118 4155 182 4219
rect 198 4155 262 4219
rect 278 4215 342 4219
rect 278 4159 282 4215
rect 282 4159 338 4215
rect 338 4159 342 4215
rect 278 4155 342 4159
rect 358 4215 422 4219
rect 358 4159 362 4215
rect 362 4159 418 4215
rect 418 4159 422 4215
rect 358 4155 422 4159
rect 438 4215 502 4219
rect 438 4159 442 4215
rect 442 4159 498 4215
rect 498 4159 502 4215
rect 438 4155 502 4159
rect 78 61 142 65
rect 78 5 82 61
rect 82 5 138 61
rect 138 5 142 61
rect 78 1 142 5
rect 158 61 222 65
rect 158 5 162 61
rect 162 5 218 61
rect 218 5 222 61
rect 158 1 222 5
rect 238 61 302 65
rect 238 5 242 61
rect 242 5 298 61
rect 298 5 302 61
rect 238 1 302 5
rect 318 61 382 65
rect 318 5 322 61
rect 322 5 378 61
rect 378 5 382 61
rect 318 1 382 5
rect 398 61 462 65
rect 398 5 402 61
rect 402 5 458 61
rect 458 5 462 61
rect 398 1 462 5
<< metal4 >>
rect 0 4219 540 4220
rect 0 4155 38 4219
rect 102 4155 118 4219
rect 182 4155 198 4219
rect 262 4155 278 4219
rect 342 4155 358 4219
rect 422 4155 438 4219
rect 502 4155 540 4219
rect 0 4154 540 4155
rect 0 126 60 4154
rect 120 66 180 4094
rect 240 126 300 4154
rect 360 66 420 4094
rect 480 126 540 4154
rect 60 65 480 66
rect 60 1 78 65
rect 142 1 158 65
rect 222 1 238 65
rect 302 1 318 65
rect 382 1 398 65
rect 462 1 480 65
rect 60 0 480 1
<< labels >>
flabel metal2 s 138 264 157 284 0 FreeSans 200 0 0 0 C0
port 1 nsew
flabel metal2 s 285 15 321 51 0 FreeSans 200 0 0 0 C1
port 2 nsew
flabel pwell s 255 566 276 615 0 FreeSans 400 0 0 0 SUB
port 3 nsew
<< properties >>
string GDS_END 29304
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 18376
string path 9.750 102.350 9.750 1.650 
string device primitive
<< end >>
