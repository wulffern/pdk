/opt/pdk/share/pdk/sky130A/libs.tech/xschem/decred_hash_macro/user_project_wrapper.spice