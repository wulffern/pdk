/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_p/end_of_life/typical/tt.spice