magic
tech sky130A
magscale 1 2
timestamp 1665766018
<< locali >>
rect 207 1548 243 1582
rect 277 1548 315 1582
rect 349 1548 387 1582
rect 421 1548 459 1582
rect 493 1548 531 1582
rect 565 1548 603 1582
rect 637 1548 675 1582
rect 709 1548 747 1582
rect 781 1548 817 1582
rect 207 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 531 54
rect 565 20 603 54
rect 637 20 675 54
rect 709 20 747 54
rect 781 20 817 54
<< viali >>
rect 243 1548 277 1582
rect 315 1548 349 1582
rect 387 1548 421 1582
rect 459 1548 493 1582
rect 531 1548 565 1582
rect 603 1548 637 1582
rect 675 1548 709 1582
rect 747 1548 781 1582
rect 243 20 277 54
rect 315 20 349 54
rect 387 20 421 54
rect 459 20 493 54
rect 531 20 565 54
rect 603 20 637 54
rect 675 20 709 54
rect 747 20 781 54
<< obsli1 >>
rect 48 1466 82 1514
rect 48 1394 82 1432
rect 48 1322 82 1360
rect 48 1250 82 1288
rect 48 1178 82 1216
rect 48 1106 82 1144
rect 48 1034 82 1072
rect 48 962 82 1000
rect 48 890 82 928
rect 48 818 82 856
rect 48 746 82 784
rect 48 674 82 712
rect 48 602 82 640
rect 48 530 82 568
rect 48 458 82 496
rect 48 386 82 424
rect 48 314 82 352
rect 48 242 82 280
rect 48 170 82 208
rect 48 88 82 136
rect 183 88 217 1514
rect 339 88 373 1514
rect 495 88 529 1514
rect 651 88 685 1514
rect 807 88 841 1514
rect 942 1466 976 1480
rect 942 1394 976 1432
rect 942 1322 976 1360
rect 942 1250 976 1288
rect 942 1178 976 1216
rect 942 1106 976 1144
rect 942 1034 976 1072
rect 942 962 976 1000
rect 942 890 976 928
rect 942 818 976 856
rect 942 746 976 784
rect 942 674 976 712
rect 942 602 976 640
rect 942 530 976 568
rect 942 458 976 496
rect 942 386 976 424
rect 942 314 976 352
rect 942 242 976 280
rect 942 170 976 208
rect 942 122 976 136
<< obsli1c >>
rect 48 1432 82 1466
rect 48 1360 82 1394
rect 48 1288 82 1322
rect 48 1216 82 1250
rect 48 1144 82 1178
rect 48 1072 82 1106
rect 48 1000 82 1034
rect 48 928 82 962
rect 48 856 82 890
rect 48 784 82 818
rect 48 712 82 746
rect 48 640 82 674
rect 48 568 82 602
rect 48 496 82 530
rect 48 424 82 458
rect 48 352 82 386
rect 48 280 82 314
rect 48 208 82 242
rect 48 136 82 170
rect 942 1432 976 1466
rect 942 1360 976 1394
rect 942 1288 976 1322
rect 942 1216 976 1250
rect 942 1144 976 1178
rect 942 1072 976 1106
rect 942 1000 976 1034
rect 942 928 976 962
rect 942 856 976 890
rect 942 784 976 818
rect 942 712 976 746
rect 942 640 976 674
rect 942 568 976 602
rect 942 496 976 530
rect 942 424 976 458
rect 942 352 976 386
rect 942 280 976 314
rect 942 208 976 242
rect 942 136 976 170
<< metal1 >>
rect 231 1582 793 1602
rect 231 1548 243 1582
rect 277 1548 315 1582
rect 349 1548 387 1582
rect 421 1548 459 1582
rect 493 1548 531 1582
rect 565 1548 603 1582
rect 637 1548 675 1582
rect 709 1548 747 1582
rect 781 1548 793 1582
rect 231 1536 793 1548
rect 36 1466 94 1497
rect 36 1432 48 1466
rect 82 1432 94 1466
rect 36 1394 94 1432
rect 36 1360 48 1394
rect 82 1360 94 1394
rect 36 1322 94 1360
rect 36 1288 48 1322
rect 82 1288 94 1322
rect 36 1250 94 1288
rect 36 1216 48 1250
rect 82 1216 94 1250
rect 36 1178 94 1216
rect 36 1144 48 1178
rect 82 1144 94 1178
rect 36 1106 94 1144
rect 36 1072 48 1106
rect 82 1072 94 1106
rect 36 1034 94 1072
rect 36 1000 48 1034
rect 82 1000 94 1034
rect 36 962 94 1000
rect 36 928 48 962
rect 82 928 94 962
rect 36 890 94 928
rect 36 856 48 890
rect 82 856 94 890
rect 36 818 94 856
rect 36 784 48 818
rect 82 784 94 818
rect 36 746 94 784
rect 36 712 48 746
rect 82 712 94 746
rect 36 674 94 712
rect 36 640 48 674
rect 82 640 94 674
rect 36 602 94 640
rect 36 568 48 602
rect 82 568 94 602
rect 36 530 94 568
rect 36 496 48 530
rect 82 496 94 530
rect 36 458 94 496
rect 36 424 48 458
rect 82 424 94 458
rect 36 386 94 424
rect 36 352 48 386
rect 82 352 94 386
rect 36 314 94 352
rect 36 280 48 314
rect 82 280 94 314
rect 36 242 94 280
rect 36 208 48 242
rect 82 208 94 242
rect 36 170 94 208
rect 36 136 48 170
rect 82 136 94 170
rect 36 105 94 136
rect 930 1466 988 1497
rect 930 1432 942 1466
rect 976 1432 988 1466
rect 930 1394 988 1432
rect 930 1360 942 1394
rect 976 1360 988 1394
rect 930 1322 988 1360
rect 930 1288 942 1322
rect 976 1288 988 1322
rect 930 1250 988 1288
rect 930 1216 942 1250
rect 976 1216 988 1250
rect 930 1178 988 1216
rect 930 1144 942 1178
rect 976 1144 988 1178
rect 930 1106 988 1144
rect 930 1072 942 1106
rect 976 1072 988 1106
rect 930 1034 988 1072
rect 930 1000 942 1034
rect 976 1000 988 1034
rect 930 962 988 1000
rect 930 928 942 962
rect 976 928 988 962
rect 930 890 988 928
rect 930 856 942 890
rect 976 856 988 890
rect 930 818 988 856
rect 930 784 942 818
rect 976 784 988 818
rect 930 746 988 784
rect 930 712 942 746
rect 976 712 988 746
rect 930 674 988 712
rect 930 640 942 674
rect 976 640 988 674
rect 930 602 988 640
rect 930 568 942 602
rect 976 568 988 602
rect 930 530 988 568
rect 930 496 942 530
rect 976 496 988 530
rect 930 458 988 496
rect 930 424 942 458
rect 976 424 988 458
rect 930 386 988 424
rect 930 352 942 386
rect 976 352 988 386
rect 930 314 988 352
rect 930 280 942 314
rect 976 280 988 314
rect 930 242 988 280
rect 930 208 942 242
rect 976 208 988 242
rect 930 170 988 208
rect 930 136 942 170
rect 976 136 988 170
rect 930 105 988 136
rect 231 54 793 66
rect 231 20 243 54
rect 277 20 315 54
rect 349 20 387 54
rect 421 20 459 54
rect 493 20 531 54
rect 565 20 603 54
rect 637 20 675 54
rect 709 20 747 54
rect 781 20 793 54
rect 231 0 793 20
<< obsm1 >>
rect 174 105 226 1497
rect 330 105 382 1497
rect 486 105 538 1497
rect 642 105 694 1497
rect 798 105 850 1497
<< metal2 >>
rect 10 1177 1014 1497
rect 10 481 1014 1121
rect 10 105 1014 425
<< labels >>
rlabel metal2 s 10 481 1014 1121 6 DRAIN
port 1 nsew
rlabel viali s 747 1548 781 1582 6 GATE
port 2 nsew
rlabel viali s 747 20 781 54 6 GATE
port 2 nsew
rlabel viali s 675 1548 709 1582 6 GATE
port 2 nsew
rlabel viali s 675 20 709 54 6 GATE
port 2 nsew
rlabel viali s 603 1548 637 1582 6 GATE
port 2 nsew
rlabel viali s 603 20 637 54 6 GATE
port 2 nsew
rlabel viali s 531 1548 565 1582 6 GATE
port 2 nsew
rlabel viali s 531 20 565 54 6 GATE
port 2 nsew
rlabel viali s 459 1548 493 1582 6 GATE
port 2 nsew
rlabel viali s 459 20 493 54 6 GATE
port 2 nsew
rlabel viali s 387 1548 421 1582 6 GATE
port 2 nsew
rlabel viali s 387 20 421 54 6 GATE
port 2 nsew
rlabel viali s 315 1548 349 1582 6 GATE
port 2 nsew
rlabel viali s 315 20 349 54 6 GATE
port 2 nsew
rlabel viali s 243 1548 277 1582 6 GATE
port 2 nsew
rlabel viali s 243 20 277 54 6 GATE
port 2 nsew
rlabel locali s 207 1548 817 1582 6 GATE
port 2 nsew
rlabel locali s 207 20 817 54 6 GATE
port 2 nsew
rlabel metal1 s 231 1536 793 1602 6 GATE
port 2 nsew
rlabel metal1 s 231 0 793 66 6 GATE
port 2 nsew
rlabel metal2 s 10 1177 1014 1497 6 SOURCE
port 3 nsew
rlabel metal2 s 10 105 1014 425 6 SOURCE
port 3 nsew
rlabel metal1 s 36 105 94 1497 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 930 105 988 1497 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 10 0 1014 1602
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4348170
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 4318450
<< end >>
