/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice