/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sky130_fd_pr__model__linear.model.spice