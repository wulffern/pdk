/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/corners/sf/specialized_cells.spice