/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/correl1.spice