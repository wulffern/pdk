magic
tech sky130B
magscale 1 2
timestamp 1665766018
<< obsli1 >>
rect 98 719 368 735
rect 98 685 108 719
rect 142 685 180 719
rect 214 685 252 719
rect 286 685 324 719
rect 358 685 368 719
rect 98 667 368 685
rect 44 605 78 621
rect 44 533 78 571
rect 44 461 78 499
rect 44 389 78 427
rect 44 317 78 355
rect 44 245 78 283
rect 44 173 78 211
rect 44 101 78 139
rect 44 51 78 67
rect 130 51 164 621
rect 216 605 250 621
rect 216 533 250 571
rect 216 461 250 499
rect 216 389 250 427
rect 216 317 250 355
rect 216 245 250 283
rect 216 173 250 211
rect 216 101 250 139
rect 216 51 250 67
rect 302 51 336 621
rect 388 605 422 621
rect 388 533 422 571
rect 388 461 422 499
rect 388 389 422 427
rect 388 317 422 355
rect 388 245 422 283
rect 388 173 422 211
rect 388 101 422 139
rect 388 51 422 67
<< obsli1c >>
rect 108 685 142 719
rect 180 685 214 719
rect 252 685 286 719
rect 324 685 358 719
rect 44 571 78 605
rect 44 499 78 533
rect 44 427 78 461
rect 44 355 78 389
rect 44 283 78 317
rect 44 211 78 245
rect 44 139 78 173
rect 44 67 78 101
rect 216 571 250 605
rect 216 499 250 533
rect 216 427 250 461
rect 216 355 250 389
rect 216 283 250 317
rect 216 211 250 245
rect 216 139 250 173
rect 216 67 250 101
rect 388 571 422 605
rect 388 499 422 533
rect 388 427 422 461
rect 388 355 422 389
rect 388 283 422 317
rect 388 211 422 245
rect 388 139 422 173
rect 388 67 422 101
<< metal1 >>
rect 96 719 370 731
rect 96 685 108 719
rect 142 685 180 719
rect 214 685 252 719
rect 286 685 324 719
rect 358 685 370 719
rect 96 673 370 685
rect 38 605 84 621
rect 38 571 44 605
rect 78 571 84 605
rect 38 533 84 571
rect 38 499 44 533
rect 78 499 84 533
rect 38 461 84 499
rect 38 427 44 461
rect 78 427 84 461
rect 38 389 84 427
rect 38 355 44 389
rect 78 355 84 389
rect 38 317 84 355
rect 38 283 44 317
rect 78 283 84 317
rect 38 245 84 283
rect 38 211 44 245
rect 78 211 84 245
rect 38 173 84 211
rect 38 139 44 173
rect 78 139 84 173
rect 38 101 84 139
rect 38 67 44 101
rect 78 67 84 101
rect 38 -29 84 67
rect 210 605 256 621
rect 210 571 216 605
rect 250 571 256 605
rect 210 533 256 571
rect 210 499 216 533
rect 250 499 256 533
rect 210 461 256 499
rect 210 427 216 461
rect 250 427 256 461
rect 210 389 256 427
rect 210 355 216 389
rect 250 355 256 389
rect 210 317 256 355
rect 210 283 216 317
rect 250 283 256 317
rect 210 245 256 283
rect 210 211 216 245
rect 250 211 256 245
rect 210 173 256 211
rect 210 139 216 173
rect 250 139 256 173
rect 210 101 256 139
rect 210 67 216 101
rect 250 67 256 101
rect 210 -29 256 67
rect 382 605 428 621
rect 382 571 388 605
rect 422 571 428 605
rect 382 533 428 571
rect 382 499 388 533
rect 422 499 428 533
rect 382 461 428 499
rect 382 427 388 461
rect 422 427 428 461
rect 382 389 428 427
rect 382 355 388 389
rect 422 355 428 389
rect 382 317 428 355
rect 382 283 388 317
rect 422 283 428 317
rect 382 245 428 283
rect 382 211 388 245
rect 422 211 428 245
rect 382 173 428 211
rect 382 139 388 173
rect 422 139 428 173
rect 382 101 428 139
rect 382 67 388 101
rect 422 67 428 101
rect 382 -29 428 67
rect 38 -89 428 -29
<< obsm1 >>
rect 121 51 173 621
rect 293 51 345 621
<< obsm2 >>
rect 114 475 180 629
rect 286 475 352 629
<< metal3 >>
rect 114 563 352 629
rect 114 475 180 563
rect 286 475 352 563
<< labels >>
rlabel metal3 s 286 475 352 563 6 DRAIN
port 1 nsew
rlabel metal3 s 114 563 352 629 6 DRAIN
port 1 nsew
rlabel metal3 s 114 475 180 563 6 DRAIN
port 1 nsew
rlabel metal1 s 96 673 370 731 6 GATE
port 2 nsew
rlabel metal1 s 382 -29 428 621 6 SOURCE
port 3 nsew
rlabel metal1 s 210 -29 256 621 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -29 84 621 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -89 428 -29 8 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 -89 466 735
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9148738
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9138218
<< end >>
