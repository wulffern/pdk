magic
tech sky130A
magscale 1 2
timestamp 1665766018
<< obsli1 >>
rect 271 2271 1996 2280
rect 271 2237 1997 2271
rect 271 2228 1996 2237
rect 93 1987 2175 2147
rect 93 325 235 1987
rect 290 1219 324 1953
rect 360 1253 394 1987
rect 430 1219 464 1953
rect 500 1253 534 1987
rect 570 1219 604 1953
rect 640 1253 674 1987
rect 710 1219 744 1953
rect 780 1253 814 1987
rect 850 1219 884 1953
rect 920 1253 954 1987
rect 990 1219 1024 1953
rect 1060 1256 1208 1987
rect 1060 1255 1180 1256
rect 290 1093 1052 1219
rect 290 359 324 1093
rect 360 325 394 1059
rect 430 359 464 1093
rect 500 325 534 1059
rect 570 359 604 1093
rect 640 325 674 1059
rect 710 359 744 1093
rect 780 325 814 1059
rect 850 359 884 1093
rect 920 325 954 1059
rect 990 359 1024 1093
rect 1088 1057 1180 1255
rect 1244 1219 1278 1953
rect 1314 1253 1348 1987
rect 1384 1219 1418 1953
rect 1454 1253 1488 1987
rect 1524 1219 1558 1953
rect 1594 1253 1628 1987
rect 1664 1219 1698 1953
rect 1734 1253 1768 1987
rect 1804 1219 1838 1953
rect 1874 1253 1908 1987
rect 1944 1219 1978 1953
rect 1216 1093 1978 1219
rect 1060 325 1208 1057
rect 1244 359 1278 1093
rect 1314 325 1348 1059
rect 1384 359 1418 1093
rect 1454 325 1488 1059
rect 1524 359 1558 1093
rect 1594 325 1628 1059
rect 1664 359 1698 1093
rect 1734 325 1768 1059
rect 1804 359 1838 1093
rect 1874 325 1908 1059
rect 1944 359 1978 1093
rect 2033 325 2175 1987
rect 93 165 2175 325
rect 271 101 1996 110
rect 271 67 1997 101
rect 271 58 1996 67
<< obsm1 >>
rect 93 2308 2175 2338
rect 93 2041 243 2308
rect 271 2071 1996 2280
rect 93 1987 1024 2041
rect 93 1897 262 1987
rect 1052 1953 1216 2071
rect 2024 2041 2175 2308
rect 1244 1987 2175 2041
rect 290 1925 1978 1953
rect 93 1869 1024 1897
rect 93 1785 262 1869
rect 1052 1841 1216 1925
rect 2006 1897 2175 1987
rect 1244 1869 2175 1897
rect 290 1813 1978 1841
rect 93 1757 1024 1785
rect 93 1673 262 1757
rect 1052 1729 1216 1813
rect 2006 1785 2175 1869
rect 1244 1757 2175 1785
rect 290 1701 1978 1729
rect 93 1645 1024 1673
rect 93 1561 262 1645
rect 1052 1617 1216 1701
rect 2006 1673 2175 1757
rect 1244 1645 2175 1673
rect 290 1589 1978 1617
rect 93 1533 1024 1561
rect 93 1449 262 1533
rect 1052 1505 1216 1589
rect 2006 1561 2175 1645
rect 1244 1533 2175 1561
rect 290 1477 1978 1505
rect 93 1421 1024 1449
rect 93 1337 262 1421
rect 1052 1393 1216 1477
rect 2006 1449 2175 1533
rect 1244 1421 2175 1449
rect 290 1365 1978 1393
rect 93 1309 1024 1337
rect 93 1003 262 1309
rect 1052 1281 1216 1365
rect 2006 1337 2175 1421
rect 1244 1309 2175 1337
rect 290 1253 1978 1281
rect 1052 1219 1216 1253
rect 290 1093 1978 1219
rect 1052 1059 1216 1093
rect 290 1031 1978 1059
rect 93 975 1024 1003
rect 93 891 262 975
rect 1052 947 1216 1031
rect 2006 1003 2175 1309
rect 1244 975 2175 1003
rect 290 919 1978 947
rect 93 863 1024 891
rect 93 779 262 863
rect 1052 835 1216 919
rect 2006 891 2175 975
rect 1244 863 2175 891
rect 290 807 1978 835
rect 93 751 1024 779
rect 93 667 262 751
rect 1052 723 1216 807
rect 2006 779 2175 863
rect 1244 751 2175 779
rect 290 695 1978 723
rect 93 639 1024 667
rect 93 555 262 639
rect 1052 611 1216 695
rect 2006 667 2175 751
rect 1244 639 2175 667
rect 290 583 1978 611
rect 93 527 1024 555
rect 93 443 262 527
rect 1052 499 1216 583
rect 2006 555 2175 639
rect 1244 527 2175 555
rect 290 471 1978 499
rect 93 415 1024 443
rect 93 325 262 415
rect 1052 387 1216 471
rect 2006 443 2175 527
rect 1244 415 2175 443
rect 290 359 1978 387
rect 93 271 1024 325
rect 93 30 243 271
rect 1052 241 1216 359
rect 2006 325 2175 415
rect 1244 271 2175 325
rect 271 58 1996 241
rect 2024 30 2175 271
rect 93 0 2175 30
<< obsm2 >>
rect 65 2071 2203 2323
rect 65 241 169 2071
rect 198 1987 1024 2041
rect 198 1953 262 1987
rect 198 1925 1024 1953
rect 198 1841 262 1925
rect 1052 1897 1216 2071
rect 1244 1987 2070 2041
rect 2006 1953 2070 1987
rect 1244 1925 2070 1953
rect 290 1869 1978 1897
rect 198 1813 1024 1841
rect 198 1729 262 1813
rect 1052 1785 1216 1869
rect 2006 1841 2070 1925
rect 1244 1813 2070 1841
rect 290 1757 1978 1785
rect 198 1701 1024 1729
rect 198 1617 262 1701
rect 1052 1673 1216 1757
rect 2006 1729 2070 1813
rect 1244 1701 2070 1729
rect 290 1645 1978 1673
rect 198 1589 1024 1617
rect 198 1505 262 1589
rect 1052 1561 1216 1645
rect 2006 1617 2070 1701
rect 1244 1589 2070 1617
rect 290 1533 1978 1561
rect 198 1477 1024 1505
rect 198 1393 262 1477
rect 1052 1449 1216 1533
rect 2006 1505 2070 1589
rect 1244 1477 2070 1505
rect 290 1421 1978 1449
rect 198 1365 1024 1393
rect 198 1281 262 1365
rect 1052 1337 1216 1421
rect 2006 1393 2070 1477
rect 1244 1365 2070 1393
rect 290 1309 1978 1337
rect 198 1253 1024 1281
rect 198 1059 262 1253
rect 1052 1219 1216 1309
rect 2006 1281 2070 1365
rect 1244 1253 2070 1281
rect 290 1093 1978 1219
rect 198 1031 1024 1059
rect 198 947 262 1031
rect 1052 1003 1216 1093
rect 2006 1059 2070 1253
rect 1244 1031 2070 1059
rect 290 975 1978 1003
rect 198 919 1024 947
rect 198 835 262 919
rect 1052 891 1216 975
rect 2006 947 2070 1031
rect 1244 919 2070 947
rect 290 863 1978 891
rect 198 807 1024 835
rect 198 723 262 807
rect 1052 779 1216 863
rect 2006 835 2070 919
rect 1244 807 2070 835
rect 290 751 1978 779
rect 198 695 1024 723
rect 198 611 262 695
rect 1052 667 1216 751
rect 2006 723 2070 807
rect 1244 695 2070 723
rect 290 639 1978 667
rect 198 583 1024 611
rect 198 499 262 583
rect 1052 555 1216 639
rect 2006 611 2070 695
rect 1244 583 2070 611
rect 290 527 1978 555
rect 198 471 1024 499
rect 198 387 262 471
rect 1052 443 1216 527
rect 2006 499 2070 583
rect 1244 471 2070 499
rect 290 415 1978 443
rect 198 359 1024 387
rect 198 325 262 359
rect 198 271 1024 325
rect 1052 241 1216 415
rect 2006 387 2070 471
rect 1244 359 2070 387
rect 2006 325 2070 359
rect 1244 271 2070 325
rect 2098 241 2203 2071
rect 65 15 2203 241
<< obsm3 >>
rect 60 15 126 2323
rect 193 2206 2075 2272
rect 193 2026 259 2206
rect 319 2086 1949 2146
rect 193 1966 1041 2026
rect 193 1786 259 1966
rect 1101 1906 1167 2086
rect 2009 2026 2075 2206
rect 1227 1966 2075 2026
rect 319 1846 1949 1906
rect 193 1726 1041 1786
rect 193 1546 259 1726
rect 1101 1666 1167 1846
rect 2009 1786 2075 1966
rect 1227 1726 2075 1786
rect 319 1606 1949 1666
rect 193 1486 1041 1546
rect 193 1306 259 1486
rect 1101 1426 1167 1606
rect 2009 1546 2075 1726
rect 1227 1486 2075 1546
rect 319 1366 1949 1426
rect 193 1246 1041 1306
rect 193 1060 259 1246
rect 1101 1186 1167 1366
rect 2009 1306 2075 1486
rect 1227 1246 2075 1306
rect 319 1120 1949 1186
rect 193 1000 1041 1060
rect 193 820 259 1000
rect 1101 940 1167 1120
rect 2009 1060 2075 1246
rect 1227 1000 2075 1060
rect 319 880 1949 940
rect 193 760 1041 820
rect 193 580 259 760
rect 1101 700 1167 880
rect 2009 820 2075 1000
rect 1227 760 2075 820
rect 319 640 1949 700
rect 193 520 1041 580
rect 193 340 259 520
rect 1101 460 1167 640
rect 2009 580 2075 760
rect 1227 520 2075 580
rect 319 400 1949 460
rect 193 280 1041 340
rect 193 100 259 280
rect 1101 220 1167 400
rect 2009 340 2075 520
rect 1227 280 2075 340
rect 319 160 1949 220
rect 2009 100 2075 280
rect 193 34 2075 100
rect 2142 15 2208 2323
<< metal4 >>
rect 60 15 126 2323
rect 193 2266 2009 2272
rect 193 2206 2075 2266
rect 193 100 259 2206
rect 319 1186 379 2146
rect 439 1246 499 2206
rect 559 1186 619 2146
rect 679 1246 739 2206
rect 799 1186 859 2146
rect 919 1246 1002 2206
rect 1062 1186 1167 2146
rect 1227 1246 1349 2206
rect 1409 1186 1469 2146
rect 1529 1246 1589 2206
rect 1649 1186 1709 2146
rect 1769 1246 1829 2206
rect 1889 1186 1949 2146
rect 319 1120 1949 1186
rect 319 160 379 1120
rect 439 100 499 1060
rect 559 160 619 1120
rect 679 100 739 1060
rect 799 160 859 1120
rect 919 100 1002 1060
rect 1062 160 1167 1120
rect 1227 100 1349 1060
rect 1409 160 1469 1120
rect 1529 100 1589 1060
rect 1649 160 1709 1120
rect 1769 100 1829 1060
rect 1889 160 1949 1120
rect 2009 100 2075 2206
rect 193 34 2075 100
rect 2142 15 2208 2323
<< metal5 >>
rect 0 0 2268 2338
<< labels >>
rlabel metal4 s 2142 15 2208 2323 6 C0
port 1 nsew
rlabel metal4 s 1889 1186 1949 2146 6 C0
port 1 nsew
rlabel metal4 s 1889 160 1949 1120 6 C0
port 1 nsew
rlabel metal4 s 1649 1186 1709 2146 6 C0
port 1 nsew
rlabel metal4 s 1649 160 1709 1120 6 C0
port 1 nsew
rlabel metal4 s 1409 1186 1469 2146 6 C0
port 1 nsew
rlabel metal4 s 1409 160 1469 1120 6 C0
port 1 nsew
rlabel metal4 s 1062 1186 1167 2146 6 C0
port 1 nsew
rlabel metal4 s 1062 160 1167 1120 6 C0
port 1 nsew
rlabel metal4 s 799 1186 859 2146 6 C0
port 1 nsew
rlabel metal4 s 799 160 859 1120 6 C0
port 1 nsew
rlabel metal4 s 559 1186 619 2146 6 C0
port 1 nsew
rlabel metal4 s 559 160 619 1120 6 C0
port 1 nsew
rlabel metal4 s 319 1186 379 2146 6 C0
port 1 nsew
rlabel metal4 s 319 1120 1949 1186 6 C0
port 1 nsew
rlabel metal4 s 319 160 379 1120 6 C0
port 1 nsew
rlabel metal4 s 60 15 126 2323 6 C0
port 1 nsew
rlabel metal4 s 2009 100 2075 2206 6 C1
port 2 nsew
rlabel metal4 s 1769 1246 1829 2206 6 C1
port 2 nsew
rlabel metal4 s 1769 100 1829 1060 6 C1
port 2 nsew
rlabel metal4 s 1529 1246 1589 2206 6 C1
port 2 nsew
rlabel metal4 s 1529 100 1589 1060 6 C1
port 2 nsew
rlabel metal4 s 1227 1246 1349 2206 6 C1
port 2 nsew
rlabel metal4 s 1227 100 1349 1060 6 C1
port 2 nsew
rlabel metal4 s 919 1246 1002 2206 6 C1
port 2 nsew
rlabel metal4 s 919 100 1002 1060 6 C1
port 2 nsew
rlabel metal4 s 679 1246 739 2206 6 C1
port 2 nsew
rlabel metal4 s 679 100 739 1060 6 C1
port 2 nsew
rlabel metal4 s 439 1246 499 2206 6 C1
port 2 nsew
rlabel metal4 s 439 100 499 1060 6 C1
port 2 nsew
rlabel metal4 s 193 2266 2009 2272 6 C1
port 2 nsew
rlabel metal4 s 193 2206 2075 2266 6 C1
port 2 nsew
rlabel metal4 s 193 100 259 2206 6 C1
port 2 nsew
rlabel metal4 s 193 34 2075 100 6 C1
port 2 nsew
rlabel metal5 s 0 0 2268 2338 6 MET5
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 2268 2338
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 702972
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 599226
string device primitive
<< end >>