/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/corners/ff/nonfet.spice