/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/lef/sky130_fd_pr.lef