magic
tech sky130A
magscale 1 2
timestamp 1665766018
<< locali >>
rect 248 1369 394 1388
rect 248 1335 262 1369
rect 296 1335 346 1369
rect 380 1335 394 1369
rect 248 1297 394 1335
rect 248 1263 262 1297
rect 296 1263 346 1297
rect 380 1263 394 1297
rect 248 1249 394 1263
rect 248 125 394 139
rect 248 91 262 125
rect 296 91 346 125
rect 380 91 394 125
rect 248 53 394 91
rect 248 19 262 53
rect 296 19 346 53
rect 380 19 394 53
rect 248 0 394 19
<< viali >>
rect 262 1335 296 1369
rect 346 1335 380 1369
rect 262 1263 296 1297
rect 346 1263 380 1297
rect 262 91 296 125
rect 346 91 380 125
rect 262 19 296 53
rect 346 19 380 53
<< obsli1 >>
rect 120 1225 186 1291
rect 456 1225 522 1291
rect 120 1203 160 1225
rect 482 1203 522 1225
rect 41 1179 160 1203
rect 41 1145 60 1179
rect 94 1145 160 1179
rect 41 1107 160 1145
rect 41 1073 60 1107
rect 94 1073 160 1107
rect 41 1035 160 1073
rect 41 1001 60 1035
rect 94 1001 160 1035
rect 41 963 160 1001
rect 41 929 60 963
rect 94 929 160 963
rect 41 891 160 929
rect 41 857 60 891
rect 94 857 160 891
rect 41 819 160 857
rect 41 785 60 819
rect 94 785 160 819
rect 41 747 160 785
rect 41 713 60 747
rect 94 713 160 747
rect 41 675 160 713
rect 41 641 60 675
rect 94 641 160 675
rect 41 603 160 641
rect 41 569 60 603
rect 94 569 160 603
rect 41 531 160 569
rect 41 497 60 531
rect 94 497 160 531
rect 41 459 160 497
rect 41 425 60 459
rect 94 425 160 459
rect 41 387 160 425
rect 41 353 60 387
rect 94 353 160 387
rect 41 315 160 353
rect 41 281 60 315
rect 94 281 160 315
rect 41 243 160 281
rect 41 209 60 243
rect 94 209 160 243
rect 41 185 160 209
rect 212 185 246 1203
rect 304 185 338 1203
rect 396 185 430 1203
rect 482 1179 601 1203
rect 482 1145 548 1179
rect 582 1145 601 1179
rect 482 1107 601 1145
rect 482 1073 548 1107
rect 582 1073 601 1107
rect 482 1035 601 1073
rect 482 1001 548 1035
rect 582 1001 601 1035
rect 482 963 601 1001
rect 482 929 548 963
rect 582 929 601 963
rect 482 891 601 929
rect 482 857 548 891
rect 582 857 601 891
rect 482 819 601 857
rect 482 785 548 819
rect 582 785 601 819
rect 482 747 601 785
rect 482 713 548 747
rect 582 713 601 747
rect 482 675 601 713
rect 482 641 548 675
rect 582 641 601 675
rect 482 603 601 641
rect 482 569 548 603
rect 582 569 601 603
rect 482 531 601 569
rect 482 497 548 531
rect 582 497 601 531
rect 482 459 601 497
rect 482 425 548 459
rect 582 425 601 459
rect 482 387 601 425
rect 482 353 548 387
rect 582 353 601 387
rect 482 315 601 353
rect 482 281 548 315
rect 582 281 601 315
rect 482 243 601 281
rect 482 209 548 243
rect 582 209 601 243
rect 482 185 601 209
rect 120 163 160 185
rect 482 163 522 185
rect 120 97 186 163
rect 456 97 522 163
<< obsli1c >>
rect 60 1145 94 1179
rect 60 1073 94 1107
rect 60 1001 94 1035
rect 60 929 94 963
rect 60 857 94 891
rect 60 785 94 819
rect 60 713 94 747
rect 60 641 94 675
rect 60 569 94 603
rect 60 497 94 531
rect 60 425 94 459
rect 60 353 94 387
rect 60 281 94 315
rect 60 209 94 243
rect 548 1145 582 1179
rect 548 1073 582 1107
rect 548 1001 582 1035
rect 548 929 582 963
rect 548 857 582 891
rect 548 785 582 819
rect 548 713 582 747
rect 548 641 582 675
rect 548 569 582 603
rect 548 497 582 531
rect 548 425 582 459
rect 548 353 582 387
rect 548 281 582 315
rect 548 209 582 243
<< metal1 >>
rect 250 1369 392 1388
rect 250 1335 262 1369
rect 296 1335 346 1369
rect 380 1335 392 1369
rect 250 1297 392 1335
rect 250 1263 262 1297
rect 296 1263 346 1297
rect 380 1263 392 1297
rect 250 1251 392 1263
rect 41 1179 100 1191
rect 41 1145 60 1179
rect 94 1145 100 1179
rect 41 1107 100 1145
rect 41 1073 60 1107
rect 94 1073 100 1107
rect 41 1035 100 1073
rect 41 1001 60 1035
rect 94 1001 100 1035
rect 41 963 100 1001
rect 41 929 60 963
rect 94 929 100 963
rect 41 891 100 929
rect 41 857 60 891
rect 94 857 100 891
rect 41 819 100 857
rect 41 785 60 819
rect 94 785 100 819
rect 41 747 100 785
rect 41 713 60 747
rect 94 713 100 747
rect 41 675 100 713
rect 41 641 60 675
rect 94 641 100 675
rect 41 603 100 641
rect 41 569 60 603
rect 94 569 100 603
rect 41 531 100 569
rect 41 497 60 531
rect 94 497 100 531
rect 41 459 100 497
rect 41 425 60 459
rect 94 425 100 459
rect 41 387 100 425
rect 41 353 60 387
rect 94 353 100 387
rect 41 315 100 353
rect 41 281 60 315
rect 94 281 100 315
rect 41 243 100 281
rect 41 209 60 243
rect 94 209 100 243
rect 41 197 100 209
rect 542 1179 601 1191
rect 542 1145 548 1179
rect 582 1145 601 1179
rect 542 1107 601 1145
rect 542 1073 548 1107
rect 582 1073 601 1107
rect 542 1035 601 1073
rect 542 1001 548 1035
rect 582 1001 601 1035
rect 542 963 601 1001
rect 542 929 548 963
rect 582 929 601 963
rect 542 891 601 929
rect 542 857 548 891
rect 582 857 601 891
rect 542 819 601 857
rect 542 785 548 819
rect 582 785 601 819
rect 542 747 601 785
rect 542 713 548 747
rect 582 713 601 747
rect 542 675 601 713
rect 542 641 548 675
rect 582 641 601 675
rect 542 603 601 641
rect 542 569 548 603
rect 582 569 601 603
rect 542 531 601 569
rect 542 497 548 531
rect 582 497 601 531
rect 542 459 601 497
rect 542 425 548 459
rect 582 425 601 459
rect 542 387 601 425
rect 542 353 548 387
rect 582 353 601 387
rect 542 315 601 353
rect 542 281 548 315
rect 582 281 601 315
rect 542 243 601 281
rect 542 209 548 243
rect 582 209 601 243
rect 542 197 601 209
rect 250 125 392 137
rect 250 91 262 125
rect 296 91 346 125
rect 380 91 392 125
rect 250 53 392 91
rect 250 19 262 53
rect 296 19 346 53
rect 380 19 392 53
rect 250 0 392 19
<< obsm1 >>
rect 203 197 255 1191
rect 295 197 347 1191
rect 387 197 439 1191
<< metal2 >>
rect 14 719 628 1191
rect 14 197 628 669
<< labels >>
rlabel metal2 s 14 719 628 1191 6 DRAIN
port 1 nsew
rlabel viali s 346 1335 380 1369 6 GATE
port 2 nsew
rlabel viali s 346 1263 380 1297 6 GATE
port 2 nsew
rlabel viali s 346 91 380 125 6 GATE
port 2 nsew
rlabel viali s 346 19 380 53 6 GATE
port 2 nsew
rlabel viali s 262 1335 296 1369 6 GATE
port 2 nsew
rlabel viali s 262 1263 296 1297 6 GATE
port 2 nsew
rlabel viali s 262 91 296 125 6 GATE
port 2 nsew
rlabel viali s 262 19 296 53 6 GATE
port 2 nsew
rlabel locali s 248 1249 394 1388 6 GATE
port 2 nsew
rlabel locali s 248 0 394 139 6 GATE
port 2 nsew
rlabel metal1 s 250 1251 392 1388 6 GATE
port 2 nsew
rlabel metal1 s 250 0 392 137 6 GATE
port 2 nsew
rlabel metal2 s 14 197 628 669 6 SOURCE
port 3 nsew
rlabel metal1 s 41 197 100 1191 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 542 197 601 1191 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 628 1388
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3783270
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3763174
string device primitive
<< end >>
