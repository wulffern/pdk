/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_e/begin_of_life/typical.spice