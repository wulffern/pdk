/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_p/begin_of_life/worst.spice