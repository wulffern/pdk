magic
tech sky130B
magscale 1 2
timestamp 1665766018
<< locali >>
rect 400 961 962 980
rect 400 855 412 961
rect 950 855 962 961
rect 400 843 962 855
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 400 0 962 19
<< viali >>
rect 412 855 950 961
rect 412 19 950 125
<< obsli1 >>
rect 190 817 256 883
rect 1106 817 1172 883
rect 190 795 230 817
rect 1132 795 1172 817
rect 41 759 230 795
rect 41 725 60 759
rect 94 725 230 759
rect 41 687 230 725
rect 41 653 60 687
rect 94 653 230 687
rect 41 615 230 653
rect 41 581 60 615
rect 94 581 230 615
rect 41 543 230 581
rect 41 509 60 543
rect 94 509 230 543
rect 41 471 230 509
rect 41 437 60 471
rect 94 437 230 471
rect 41 399 230 437
rect 41 365 60 399
rect 94 365 230 399
rect 41 327 230 365
rect 41 293 60 327
rect 94 293 230 327
rect 41 255 230 293
rect 41 221 60 255
rect 94 221 230 255
rect 41 185 230 221
rect 352 185 386 795
rect 508 185 542 795
rect 664 185 698 795
rect 820 185 854 795
rect 976 185 1010 795
rect 1132 759 1321 795
rect 1132 725 1268 759
rect 1302 725 1321 759
rect 1132 687 1321 725
rect 1132 653 1268 687
rect 1302 653 1321 687
rect 1132 615 1321 653
rect 1132 581 1268 615
rect 1302 581 1321 615
rect 1132 543 1321 581
rect 1132 509 1268 543
rect 1302 509 1321 543
rect 1132 471 1321 509
rect 1132 437 1268 471
rect 1302 437 1321 471
rect 1132 399 1321 437
rect 1132 365 1268 399
rect 1302 365 1321 399
rect 1132 327 1321 365
rect 1132 293 1268 327
rect 1302 293 1321 327
rect 1132 255 1321 293
rect 1132 221 1268 255
rect 1302 221 1321 255
rect 1132 185 1321 221
rect 190 163 230 185
rect 1132 163 1172 185
rect 190 97 256 163
rect 1106 97 1172 163
<< obsli1c >>
rect 60 725 94 759
rect 60 653 94 687
rect 60 581 94 615
rect 60 509 94 543
rect 60 437 94 471
rect 60 365 94 399
rect 60 293 94 327
rect 60 221 94 255
rect 1268 725 1302 759
rect 1268 653 1302 687
rect 1268 581 1302 615
rect 1268 509 1302 543
rect 1268 437 1302 471
rect 1268 365 1302 399
rect 1268 293 1302 327
rect 1268 221 1302 255
<< metal1 >>
rect 400 961 962 980
rect 400 855 412 961
rect 950 855 962 961
rect 400 843 962 855
rect 41 759 100 771
rect 41 725 60 759
rect 94 725 100 759
rect 41 687 100 725
rect 41 653 60 687
rect 94 653 100 687
rect 41 615 100 653
rect 41 581 60 615
rect 94 581 100 615
rect 41 543 100 581
rect 41 509 60 543
rect 94 509 100 543
rect 41 471 100 509
rect 41 437 60 471
rect 94 437 100 471
rect 41 399 100 437
rect 41 365 60 399
rect 94 365 100 399
rect 41 327 100 365
rect 41 293 60 327
rect 94 293 100 327
rect 41 255 100 293
rect 41 221 60 255
rect 94 221 100 255
rect 41 209 100 221
rect 1262 759 1321 771
rect 1262 725 1268 759
rect 1302 725 1321 759
rect 1262 687 1321 725
rect 1262 653 1268 687
rect 1302 653 1321 687
rect 1262 615 1321 653
rect 1262 581 1268 615
rect 1302 581 1321 615
rect 1262 543 1321 581
rect 1262 509 1268 543
rect 1302 509 1321 543
rect 1262 471 1321 509
rect 1262 437 1268 471
rect 1302 437 1321 471
rect 1262 399 1321 437
rect 1262 365 1268 399
rect 1302 365 1321 399
rect 1262 327 1321 365
rect 1262 293 1268 327
rect 1302 293 1321 327
rect 1262 255 1321 293
rect 1262 221 1268 255
rect 1302 221 1321 255
rect 1262 209 1321 221
rect 400 125 962 137
rect 400 19 412 125
rect 950 19 962 125
rect 400 0 962 19
<< obsm1 >>
rect 343 209 395 771
rect 499 209 551 771
rect 655 209 707 771
rect 811 209 863 771
rect 967 209 1019 771
<< metal2 >>
rect 14 515 1348 771
rect 14 209 1348 465
<< labels >>
rlabel metal2 s 14 515 1348 771 6 DRAIN
port 1 nsew
rlabel viali s 412 855 950 961 6 GATE
port 2 nsew
rlabel viali s 412 19 950 125 6 GATE
port 2 nsew
rlabel locali s 400 843 962 980 6 GATE
port 2 nsew
rlabel locali s 400 0 962 137 6 GATE
port 2 nsew
rlabel metal1 s 400 843 962 980 6 GATE
port 2 nsew
rlabel metal1 s 400 0 962 137 6 GATE
port 2 nsew
rlabel metal2 s 14 209 1348 465 6 SOURCE
port 3 nsew
rlabel metal1 s 41 209 100 771 6 SUBSTRATE
port 4 nsew
rlabel metal1 s 1262 209 1321 771 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 14 0 1348 980
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 8485672
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 8463118
string device primitive
<< end >>
