/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_see/begin_of_life/worst.spice