/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_see_p/end_of_life/ff.spice