/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/correl3.spice