magic
tech sky130B
magscale 1 2
timestamp 1665766018
<< locali >>
rect 217 1160 255 1194
rect 289 1160 327 1194
rect 361 1160 399 1194
rect 433 1160 471 1194
rect 505 1160 543 1194
rect 577 1160 615 1194
rect 649 1160 687 1194
rect 721 1160 759 1194
rect 48 1020 82 1058
rect 48 948 82 986
rect 48 876 82 914
rect 48 804 82 842
rect 48 732 82 770
rect 48 660 82 698
rect 48 588 82 626
rect 48 516 82 554
rect 48 444 82 482
rect 48 372 82 410
rect 48 300 82 338
rect 48 228 82 266
rect 48 122 82 194
rect 894 1020 928 1058
rect 894 948 928 986
rect 894 876 928 914
rect 894 804 928 842
rect 894 732 928 770
rect 894 660 928 698
rect 894 588 928 626
rect 894 516 928 554
rect 894 444 928 482
rect 894 372 928 410
rect 894 300 928 338
rect 894 228 928 266
rect 894 122 928 194
rect 217 20 255 54
rect 289 20 327 54
rect 361 20 399 54
rect 433 20 471 54
rect 505 20 543 54
rect 577 20 615 54
rect 649 20 687 54
rect 721 20 759 54
<< viali >>
rect 183 1160 217 1194
rect 255 1160 289 1194
rect 327 1160 361 1194
rect 399 1160 433 1194
rect 471 1160 505 1194
rect 543 1160 577 1194
rect 615 1160 649 1194
rect 687 1160 721 1194
rect 759 1160 793 1194
rect 48 1058 82 1092
rect 48 986 82 1020
rect 48 914 82 948
rect 48 842 82 876
rect 48 770 82 804
rect 48 698 82 732
rect 48 626 82 660
rect 48 554 82 588
rect 48 482 82 516
rect 48 410 82 444
rect 48 338 82 372
rect 48 266 82 300
rect 48 194 82 228
rect 894 1058 928 1092
rect 894 986 928 1020
rect 894 914 928 948
rect 894 842 928 876
rect 894 770 928 804
rect 894 698 928 732
rect 894 626 928 660
rect 894 554 928 588
rect 894 482 928 516
rect 894 410 928 444
rect 894 338 928 372
rect 894 266 928 300
rect 894 194 928 228
rect 183 20 217 54
rect 255 20 289 54
rect 327 20 361 54
rect 399 20 433 54
rect 471 20 505 54
rect 543 20 577 54
rect 615 20 649 54
rect 687 20 721 54
rect 759 20 793 54
<< obsli1 >>
rect 159 98 193 1116
rect 315 98 349 1116
rect 471 98 505 1116
rect 627 98 661 1116
rect 783 98 817 1116
<< metal1 >>
rect 171 1194 805 1214
rect 171 1160 183 1194
rect 217 1160 255 1194
rect 289 1160 327 1194
rect 361 1160 399 1194
rect 433 1160 471 1194
rect 505 1160 543 1194
rect 577 1160 615 1194
rect 649 1160 687 1194
rect 721 1160 759 1194
rect 793 1160 805 1194
rect 171 1148 805 1160
rect 36 1092 94 1104
rect 36 1058 48 1092
rect 82 1058 94 1092
rect 36 1020 94 1058
rect 36 986 48 1020
rect 82 986 94 1020
rect 36 948 94 986
rect 36 914 48 948
rect 82 914 94 948
rect 36 876 94 914
rect 36 842 48 876
rect 82 842 94 876
rect 36 804 94 842
rect 36 770 48 804
rect 82 770 94 804
rect 36 732 94 770
rect 36 698 48 732
rect 82 698 94 732
rect 36 660 94 698
rect 36 626 48 660
rect 82 626 94 660
rect 36 588 94 626
rect 36 554 48 588
rect 82 554 94 588
rect 36 516 94 554
rect 36 482 48 516
rect 82 482 94 516
rect 36 444 94 482
rect 36 410 48 444
rect 82 410 94 444
rect 36 372 94 410
rect 36 338 48 372
rect 82 338 94 372
rect 36 300 94 338
rect 36 266 48 300
rect 82 266 94 300
rect 36 228 94 266
rect 36 194 48 228
rect 82 194 94 228
rect 36 110 94 194
rect 882 1092 940 1104
rect 882 1058 894 1092
rect 928 1058 940 1092
rect 882 1020 940 1058
rect 882 986 894 1020
rect 928 986 940 1020
rect 882 948 940 986
rect 882 914 894 948
rect 928 914 940 948
rect 882 876 940 914
rect 882 842 894 876
rect 928 842 940 876
rect 882 804 940 842
rect 882 770 894 804
rect 928 770 940 804
rect 882 732 940 770
rect 882 698 894 732
rect 928 698 940 732
rect 882 660 940 698
rect 882 626 894 660
rect 928 626 940 660
rect 882 588 940 626
rect 882 554 894 588
rect 928 554 940 588
rect 882 516 940 554
rect 882 482 894 516
rect 928 482 940 516
rect 882 444 940 482
rect 882 410 894 444
rect 928 410 940 444
rect 882 372 940 410
rect 882 338 894 372
rect 928 338 940 372
rect 882 300 940 338
rect 882 266 894 300
rect 928 266 940 300
rect 882 228 940 266
rect 882 194 894 228
rect 928 194 940 228
rect 882 110 940 194
rect 171 54 805 66
rect 171 20 183 54
rect 217 20 255 54
rect 289 20 327 54
rect 361 20 399 54
rect 433 20 471 54
rect 505 20 543 54
rect 577 20 615 54
rect 649 20 687 54
rect 721 20 759 54
rect 793 20 805 54
rect 171 0 805 20
<< obsm1 >>
rect 150 110 202 1104
rect 306 110 358 1104
rect 462 110 514 1104
rect 618 110 670 1104
rect 774 110 826 1104
<< metal2 >>
rect 10 632 966 1104
rect 10 110 966 582
<< labels >>
rlabel viali s 894 1058 928 1092 6 BULK
port 1 nsew
rlabel viali s 894 986 928 1020 6 BULK
port 1 nsew
rlabel viali s 894 914 928 948 6 BULK
port 1 nsew
rlabel viali s 894 842 928 876 6 BULK
port 1 nsew
rlabel viali s 894 770 928 804 6 BULK
port 1 nsew
rlabel viali s 894 698 928 732 6 BULK
port 1 nsew
rlabel viali s 894 626 928 660 6 BULK
port 1 nsew
rlabel viali s 894 554 928 588 6 BULK
port 1 nsew
rlabel viali s 894 482 928 516 6 BULK
port 1 nsew
rlabel viali s 894 410 928 444 6 BULK
port 1 nsew
rlabel viali s 894 338 928 372 6 BULK
port 1 nsew
rlabel viali s 894 266 928 300 6 BULK
port 1 nsew
rlabel viali s 894 194 928 228 6 BULK
port 1 nsew
rlabel viali s 48 1058 82 1092 6 BULK
port 1 nsew
rlabel viali s 48 986 82 1020 6 BULK
port 1 nsew
rlabel viali s 48 914 82 948 6 BULK
port 1 nsew
rlabel viali s 48 842 82 876 6 BULK
port 1 nsew
rlabel viali s 48 770 82 804 6 BULK
port 1 nsew
rlabel viali s 48 698 82 732 6 BULK
port 1 nsew
rlabel viali s 48 626 82 660 6 BULK
port 1 nsew
rlabel viali s 48 554 82 588 6 BULK
port 1 nsew
rlabel viali s 48 482 82 516 6 BULK
port 1 nsew
rlabel viali s 48 410 82 444 6 BULK
port 1 nsew
rlabel viali s 48 338 82 372 6 BULK
port 1 nsew
rlabel viali s 48 266 82 300 6 BULK
port 1 nsew
rlabel viali s 48 194 82 228 6 BULK
port 1 nsew
rlabel locali s 894 122 928 1092 6 BULK
port 1 nsew
rlabel locali s 48 122 82 1092 6 BULK
port 1 nsew
rlabel metal1 s 882 110 940 1104 6 BULK
port 1 nsew
rlabel metal1 s 36 110 94 1104 6 BULK
port 1 nsew
rlabel metal2 s 10 632 966 1104 6 DRAIN
port 2 nsew
rlabel viali s 759 1160 793 1194 6 GATE
port 3 nsew
rlabel viali s 759 20 793 54 6 GATE
port 3 nsew
rlabel viali s 687 1160 721 1194 6 GATE
port 3 nsew
rlabel viali s 687 20 721 54 6 GATE
port 3 nsew
rlabel viali s 615 1160 649 1194 6 GATE
port 3 nsew
rlabel viali s 615 20 649 54 6 GATE
port 3 nsew
rlabel viali s 543 1160 577 1194 6 GATE
port 3 nsew
rlabel viali s 543 20 577 54 6 GATE
port 3 nsew
rlabel viali s 471 1160 505 1194 6 GATE
port 3 nsew
rlabel viali s 471 20 505 54 6 GATE
port 3 nsew
rlabel viali s 399 1160 433 1194 6 GATE
port 3 nsew
rlabel viali s 399 20 433 54 6 GATE
port 3 nsew
rlabel viali s 327 1160 361 1194 6 GATE
port 3 nsew
rlabel viali s 327 20 361 54 6 GATE
port 3 nsew
rlabel viali s 255 1160 289 1194 6 GATE
port 3 nsew
rlabel viali s 255 20 289 54 6 GATE
port 3 nsew
rlabel viali s 183 1160 217 1194 6 GATE
port 3 nsew
rlabel viali s 183 20 217 54 6 GATE
port 3 nsew
rlabel locali s 183 1160 793 1194 6 GATE
port 3 nsew
rlabel locali s 183 20 793 54 6 GATE
port 3 nsew
rlabel metal1 s 171 1148 805 1214 6 GATE
port 3 nsew
rlabel metal1 s 171 0 805 66 6 GATE
port 3 nsew
rlabel metal2 s 10 110 966 582 6 SOURCE
port 4 nsew
<< properties >>
string FIXED_BBOX 0 0 976 1214
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 10051678
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10029198
<< end >>
