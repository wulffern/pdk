/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/corners/leak/rf.spice