magic
tech sky130B
magscale 1 2
timestamp 1665766018
<< obsli1 >>
rect 98 519 368 535
rect 98 485 108 519
rect 142 485 180 519
rect 214 485 252 519
rect 286 485 324 519
rect 358 485 368 519
rect 98 467 368 485
rect 44 397 78 421
rect 44 325 78 363
rect 44 253 78 291
rect 44 181 78 219
rect 44 109 78 147
rect 44 51 78 75
rect 130 51 164 421
rect 216 397 250 421
rect 216 325 250 363
rect 216 253 250 291
rect 216 181 250 219
rect 216 109 250 147
rect 216 51 250 75
rect 302 51 336 421
rect 388 397 422 421
rect 388 325 422 363
rect 388 253 422 291
rect 388 181 422 219
rect 388 109 422 147
rect 388 51 422 75
<< obsli1c >>
rect 108 485 142 519
rect 180 485 214 519
rect 252 485 286 519
rect 324 485 358 519
rect 44 363 78 397
rect 44 291 78 325
rect 44 219 78 253
rect 44 147 78 181
rect 44 75 78 109
rect 216 363 250 397
rect 216 291 250 325
rect 216 219 250 253
rect 216 147 250 181
rect 216 75 250 109
rect 388 363 422 397
rect 388 291 422 325
rect 388 219 422 253
rect 388 147 422 181
rect 388 75 422 109
<< metal1 >>
rect 96 519 370 531
rect 96 485 108 519
rect 142 485 180 519
rect 214 485 252 519
rect 286 485 324 519
rect 358 485 370 519
rect 96 473 370 485
rect 38 397 84 421
rect 38 363 44 397
rect 78 363 84 397
rect 38 325 84 363
rect 38 291 44 325
rect 78 291 84 325
rect 38 253 84 291
rect 38 219 44 253
rect 78 219 84 253
rect 38 181 84 219
rect 38 147 44 181
rect 78 147 84 181
rect 38 109 84 147
rect 38 75 44 109
rect 78 75 84 109
rect 38 -29 84 75
rect 210 397 256 421
rect 210 363 216 397
rect 250 363 256 397
rect 210 325 256 363
rect 210 291 216 325
rect 250 291 256 325
rect 210 253 256 291
rect 210 219 216 253
rect 250 219 256 253
rect 210 181 256 219
rect 210 147 216 181
rect 250 147 256 181
rect 210 109 256 147
rect 210 75 216 109
rect 250 75 256 109
rect 210 -29 256 75
rect 382 397 428 421
rect 382 363 388 397
rect 422 363 428 397
rect 382 325 428 363
rect 382 291 388 325
rect 422 291 428 325
rect 382 253 428 291
rect 382 219 388 253
rect 422 219 428 253
rect 382 181 428 219
rect 382 147 388 181
rect 422 147 428 181
rect 382 109 428 147
rect 382 75 388 109
rect 422 75 428 109
rect 382 -29 428 75
rect 38 -89 428 -29
<< obsm1 >>
rect 121 51 173 421
rect 293 51 345 421
<< obsm2 >>
rect 114 275 180 429
rect 286 275 352 429
<< metal3 >>
rect 114 363 352 429
rect 114 275 180 363
rect 286 275 352 363
<< labels >>
rlabel metal3 s 286 275 352 363 6 DRAIN
port 1 nsew
rlabel metal3 s 114 363 352 429 6 DRAIN
port 1 nsew
rlabel metal3 s 114 275 180 363 6 DRAIN
port 1 nsew
rlabel metal1 s 96 473 370 531 6 GATE
port 2 nsew
rlabel metal1 s 382 -29 428 421 6 SOURCE
port 3 nsew
rlabel metal1 s 210 -29 256 421 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -29 84 421 6 SOURCE
port 3 nsew
rlabel metal1 s 38 -89 428 -29 8 SOURCE
port 3 nsew
<< properties >>
string FIXED_BBOX 0 -89 466 535
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 9138144
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 9129544
<< end >>
