/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/parameters/fast_70p.spice