/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_see_e/end_of_life/typical.spice