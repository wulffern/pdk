/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos_e/end_of_life/ff.spice