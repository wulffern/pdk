magic
tech sky130B
magscale 1 2
timestamp 1665766018
<< pwell >>
rect 74 370 90 389
<< obsli1 >>
rect 101 447 371 463
rect 101 413 111 447
rect 145 413 183 447
rect 217 413 255 447
rect 289 413 327 447
rect 361 413 371 447
rect 101 397 371 413
rect 47 329 81 357
rect 47 257 81 295
rect 47 185 81 223
rect 47 113 81 151
rect 47 51 81 79
rect 133 51 167 357
rect 219 329 253 357
rect 219 257 253 295
rect 219 185 253 223
rect 219 113 253 151
rect 219 51 253 79
rect 305 51 339 357
rect 391 329 425 357
rect 391 257 425 295
rect 391 185 425 223
rect 391 113 425 151
rect 391 51 425 79
<< obsli1c >>
rect 111 413 145 447
rect 183 413 217 447
rect 255 413 289 447
rect 327 413 361 447
rect 47 295 81 329
rect 47 223 81 257
rect 47 151 81 185
rect 47 79 81 113
rect 219 295 253 329
rect 219 223 253 257
rect 219 151 253 185
rect 219 79 253 113
rect 391 295 425 329
rect 391 223 425 257
rect 391 151 425 185
rect 391 79 425 113
<< metal1 >>
rect 99 447 373 459
rect 99 413 111 447
rect 145 413 183 447
rect 217 413 255 447
rect 289 413 327 447
rect 361 413 373 447
rect 99 401 373 413
rect 41 329 87 357
rect 41 295 47 329
rect 81 295 87 329
rect 41 257 87 295
rect 41 223 47 257
rect 81 223 87 257
rect 41 185 87 223
rect 41 151 47 185
rect 81 151 87 185
rect 41 113 87 151
rect 41 79 47 113
rect 81 79 87 113
rect 41 -29 87 79
rect 213 329 259 357
rect 213 295 219 329
rect 253 295 259 329
rect 213 257 259 295
rect 213 223 219 257
rect 253 223 259 257
rect 213 185 259 223
rect 213 151 219 185
rect 253 151 259 185
rect 213 113 259 151
rect 213 79 219 113
rect 253 79 259 113
rect 213 -29 259 79
rect 385 329 431 357
rect 385 295 391 329
rect 425 295 431 329
rect 385 257 431 295
rect 385 223 391 257
rect 425 223 431 257
rect 385 185 431 223
rect 385 151 391 185
rect 425 151 431 185
rect 385 113 431 151
rect 385 79 391 113
rect 425 79 431 113
rect 385 -29 431 79
rect 41 -89 431 -29
<< obsm1 >>
rect 124 51 176 357
rect 296 51 348 357
<< obsm2 >>
rect 117 203 183 357
rect 289 203 355 357
<< metal3 >>
rect 117 291 355 357
rect 117 203 183 291
rect 289 203 355 291
<< labels >>
rlabel metal3 s 289 203 355 291 6 DRAIN
port 1 nsew
rlabel metal3 s 117 291 355 357 6 DRAIN
port 1 nsew
rlabel metal3 s 117 203 183 291 6 DRAIN
port 1 nsew
rlabel metal1 s 99 401 373 459 6 GATE
port 2 nsew
rlabel metal1 s 385 -29 431 357 6 SOURCE
port 3 nsew
rlabel metal1 s 213 -29 259 357 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -29 87 357 6 SOURCE
port 3 nsew
rlabel metal1 s 41 -89 431 -29 8 SOURCE
port 3 nsew
rlabel pwell s 74 370 90 389 6 SUBSTRATE
port 4 nsew
<< properties >>
string FIXED_BBOX 36 -89 436 463
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 3327492
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 3319526
<< end >>
