/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/r+c.mrp1monte.spice