/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__nfet_20v0_reverse_iso__subcircuit.pm3.spice