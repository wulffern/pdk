/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/parameters/critical.spice