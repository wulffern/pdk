/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/correl2.spice