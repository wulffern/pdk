/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos/begin_of_life/typical.spice