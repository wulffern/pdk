/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/corners/ff/specialized_cells.spice