magic
tech sky130B
magscale 1 2
timestamp 1665766018
<< obsm2 >>
rect -4079 11002 -689 12502
tri -689 11002 811 12502 sw
tri -1311 9000 691 11002 ne
rect 691 10500 811 11002
tri 811 10500 1313 11002 sw
rect 691 9000 4024 10500
rect 6408 -750 15500 750
tri -1311 -13004 691 -11002 se
rect 691 -12502 3925 -11002
rect 691 -13004 811 -12502
tri 811 -13004 1313 -12502 nw
rect -4123 -14504 -689 -13004
tri -689 -14504 811 -13004 nw
<< obsm3 >>
tri -7509 13004 -6009 14504 se
rect -6009 13004 6009 14504
tri -9136 11377 -7509 13004 se
rect -7509 12375 -6016 13004
tri -6016 12375 -5387 13004 nw
tri 5387 12502 5889 13004 ne
rect 5889 12502 6009 13004
tri 6009 12502 8011 14504 sw
tri -5307 12375 -5180 12502 se
rect -5180 12375 -1739 12502
rect -7509 11871 -6520 12375
tri -6520 11871 -6016 12375 nw
tri -5811 11871 -5307 12375 se
rect -5307 12228 -1739 12375
tri -1739 12228 -1465 12502 sw
rect -5307 11871 -1453 12228
rect -7509 11377 -7014 11871
tri -7014 11377 -6520 11871 nw
tri -6305 11377 -5811 11871 se
rect -5811 11377 -1453 11871
tri -10883 9630 -9136 11377 se
rect -9136 11089 -7302 11377
tri -7302 11089 -7014 11377 nw
tri -6593 11089 -6305 11377 se
rect -6305 11276 -1453 11377
rect -6305 11089 -1739 11276
rect -9136 10380 -8011 11089
tri -8011 10380 -7302 11089 nw
tri -7302 10380 -6593 11089 se
rect -6593 11002 -1739 11089
tri -1739 11002 -1465 11276 nw
rect -6593 10380 -5180 11002
tri -5180 10380 -4558 11002 nw
tri -1313 10500 689 12502 se
rect 689 12255 5180 12502
tri 5180 12255 5427 12502 sw
tri 5889 12255 6136 12502 ne
rect 6136 12375 8011 12502
tri 8011 12375 8138 12502 sw
rect 6136 12255 8138 12375
tri 8138 12255 8258 12375 sw
rect 689 11546 5427 12255
tri 5427 11546 6136 12255 sw
tri 6136 11546 6845 12255 ne
rect 6845 11546 8258 12255
rect 689 11002 6136 11546
rect 689 10500 809 11002
tri 809 10500 1311 11002 nw
tri 4558 10500 5060 11002 ne
rect 5060 10837 6136 11002
tri 6136 10837 6845 11546 sw
tri 6845 10837 7554 11546 ne
rect 7554 10837 8258 11546
rect 5060 10500 6845 10837
tri -4471 10380 -4351 10500 se
rect -4351 10380 689 10500
tri 689 10380 809 10500 nw
rect -9136 9868 -8523 10380
tri -8523 9868 -8011 10380 nw
tri -7814 9868 -7302 10380 se
rect -7302 9868 -5692 10380
tri -5692 9868 -5180 10380 nw
tri -4983 9868 -4471 10380 se
rect -4471 9868 -691 10380
rect -9136 9630 -8761 9868
tri -8761 9630 -8523 9868 nw
tri -8052 9630 -7814 9868 se
rect -7814 9630 -6186 9868
tri -12382 8131 -10883 9630 se
rect -10883 8967 -9424 9630
tri -9424 8967 -8761 9630 nw
tri -8715 8967 -8052 9630 se
rect -8052 9374 -6186 9630
tri -6186 9374 -5692 9868 nw
tri -5477 9374 -4983 9868 se
rect -4983 9374 -691 9868
rect -8052 8967 -6593 9374
tri -6593 8967 -6186 9374 nw
tri -5884 8967 -5477 9374 se
rect -5477 9000 -691 9374
tri -691 9000 689 10380 nw
tri 1410 10226 1684 10500 se
rect 1684 10253 4351 10500
tri 4351 10253 4598 10500 sw
tri 5060 10253 5307 10500 ne
rect 5307 10253 6845 10500
rect 1684 10226 4598 10253
rect 1410 9671 4598 10226
tri 4598 9671 5180 10253 sw
tri 5307 9671 5889 10253 ne
rect 5889 10133 6845 10253
tri 6845 10133 7549 10837 sw
tri 7554 10133 8258 10837 ne
tri 8258 10133 10380 12255 sw
rect 5889 9671 7549 10133
rect 1410 9274 5180 9671
tri 1410 9000 1684 9274 ne
rect 1684 9000 5180 9274
tri 5180 9000 5851 9671 sw
tri 5889 9000 6560 9671 ne
rect 6560 9424 7549 9671
tri 7549 9424 8258 10133 sw
tri 8258 9424 8967 10133 ne
rect 8967 9424 10380 10133
rect 6560 9000 8258 9424
rect -5477 8967 -5307 9000
rect -10883 8258 -10133 8967
tri -10133 8258 -9424 8967 nw
tri -9424 8258 -8715 8967 se
rect -8715 8258 -7302 8967
tri -7302 8258 -6593 8967 nw
tri -6593 8258 -5884 8967 se
rect -5884 8258 -5307 8967
rect -10883 8131 -10260 8258
tri -10260 8131 -10133 8258 nw
tri -9551 8131 -9424 8258 se
rect -9424 8131 -7429 8258
tri -7429 8131 -7302 8258 nw
tri -6720 8131 -6593 8258 se
rect -6593 8131 -5307 8258
tri -14504 6009 -12382 8131 se
rect -12382 7422 -10969 8131
tri -10969 7422 -10260 8131 nw
tri -10260 7422 -9551 8131 se
rect -9551 7422 -8138 8131
tri -8138 7422 -7429 8131 nw
tri -7429 7422 -6720 8131 se
rect -6720 7422 -5307 8131
tri -5307 7422 -3729 9000 nw
rect -12382 6845 -11546 7422
tri -11546 6845 -10969 7422 nw
tri -10837 6845 -10260 7422 se
rect -10260 6845 -8715 7422
tri -8715 6845 -8138 7422 nw
tri -8006 6845 -7429 7422 se
rect -7429 6845 -6720 7422
rect -12382 6136 -12255 6845
tri -12255 6136 -11546 6845 nw
tri -11546 6136 -10837 6845 se
rect -10837 6136 -9424 6845
tri -9424 6136 -8715 6845 nw
tri -8715 6136 -8006 6845 se
rect -8006 6136 -6720 6845
tri -12382 6009 -12255 6136 nw
tri -11673 6009 -11546 6136 se
rect -11546 6009 -9671 6136
rect -14504 -6009 -13004 6009
tri -13004 5387 -12382 6009 nw
tri -12295 5387 -11673 6009 se
rect -11673 5889 -9671 6009
tri -9671 5889 -9424 6136 nw
tri -8962 5889 -8715 6136 se
rect -8715 6009 -6720 6136
tri -6720 6009 -5307 7422 nw
tri 3729 6965 5764 9000 ne
rect 5764 8595 5851 9000
tri 5851 8595 6256 9000 sw
tri 6560 8595 6965 9000 ne
rect 6965 8715 8258 9000
tri 8258 8715 8967 9424 sw
tri 8967 9000 9391 9424 ne
rect 9391 9000 10380 9424
tri 9391 8715 9676 9000 ne
rect 9676 8715 10380 9000
rect 6965 8595 8967 8715
rect 5764 8131 6256 8595
tri 6256 8131 6720 8595 sw
tri 6965 8131 7429 8595 ne
rect 7429 8131 8967 8595
rect 5764 7422 6720 8131
tri 6720 7422 7429 8131 sw
tri 7429 7422 8138 8131 ne
rect 8138 8011 8967 8131
tri 8967 8011 9671 8715 sw
tri 9676 8011 10380 8715 ne
tri 10380 8011 12502 10133 sw
rect 8138 7422 9671 8011
rect 5764 7182 7429 7422
tri 7429 7182 7669 7422 sw
tri 8138 7302 8258 7422 ne
rect 8258 7302 9671 7422
tri 9671 7302 10380 8011 sw
tri 10380 7302 11089 8011 ne
rect 11089 7302 12502 8011
tri 8258 7182 8378 7302 ne
rect 8378 7182 10380 7302
rect 5764 6965 7669 7182
tri 5764 6256 6473 6965 ne
rect 6473 6473 7669 6965
tri 7669 6473 8378 7182 sw
tri 8378 6473 9087 7182 ne
rect 9087 6593 10380 7182
tri 10380 6593 11089 7302 sw
tri 11089 7182 11209 7302 ne
rect 11209 7182 12502 7302
tri 11209 6593 11798 7182 ne
rect 11798 6593 12502 7182
rect 9087 6473 11089 6593
rect 6473 6256 8378 6473
tri 6473 6009 6720 6256 ne
rect 6720 6009 8378 6256
tri 8378 6009 8842 6473 sw
tri 9087 6009 9551 6473 ne
rect 9551 6009 11089 6473
rect -8715 5889 -8378 6009
rect -11673 5387 -10380 5889
tri -12502 5180 -12295 5387 se
rect -12295 5180 -10380 5387
tri -10380 5180 -9671 5889 nw
tri -9671 5180 -8962 5889 se
rect -8962 5180 -8378 5889
rect -12502 -5180 -11002 5180
tri -11002 4558 -10380 5180 nw
tri -10293 4558 -9671 5180 se
rect -9671 4558 -8378 5180
tri -10500 4351 -10293 4558 se
rect -10293 4351 -8378 4558
tri -8378 4351 -6720 6009 nw
tri 6720 4351 8378 6009 ne
rect 8378 5387 8842 6009
tri 8842 5387 9464 6009 sw
tri 9551 5387 10173 6009 ne
rect 10173 5889 11089 6009
tri 11089 5889 11793 6593 sw
tri 11798 5889 12502 6593 ne
tri 12502 6009 14504 8011 sw
rect 12502 5889 14504 6009
rect 10173 5387 11793 5889
rect 8378 5060 9464 5387
tri 9464 5060 9791 5387 sw
tri 10173 5060 10500 5387 ne
rect 10500 5180 11793 5387
tri 11793 5180 12502 5889 sw
tri 12502 5387 13004 5889 ne
rect 10500 5060 12502 5180
rect 8378 4351 9791 5060
tri 9791 4351 10500 5060 sw
tri 10500 4558 11002 5060 ne
rect -10500 750 -9000 4351
tri -9000 3729 -8378 4351 nw
tri 8378 3729 9000 4351 ne
rect -10500 -750 8000 750
rect -10500 -4351 -9000 -750
tri -10500 -4558 -10293 -4351 ne
rect -10293 -4558 -9000 -4351
tri -11002 -5180 -10380 -4558 sw
tri -10293 -5180 -9671 -4558 ne
rect -9671 -5180 -9000 -4558
tri -12502 -5387 -12295 -5180 ne
rect -12295 -5387 -10380 -5180
tri -13004 -6009 -12382 -5387 sw
tri -12295 -5889 -11793 -5387 ne
rect -11793 -5889 -10380 -5387
tri -10380 -5889 -9671 -5180 sw
tri -9671 -5387 -9464 -5180 ne
rect -9464 -5387 -9000 -5180
tri -9000 -5387 -7342 -3729 sw
tri 7342 -5387 9000 -3729 se
rect 9000 -4351 10500 4351
rect 9000 -5060 9791 -4351
tri 9791 -5060 10500 -4351 nw
tri 10500 -5060 11002 -4558 se
rect 11002 -5060 12502 5060
rect 13004 3250 14504 5889
rect 13004 1750 15500 3250
rect 9000 -5387 9464 -5060
tri 9464 -5387 9791 -5060 nw
tri 10173 -5387 10500 -5060 se
rect 10500 -5180 12502 -5060
rect 10500 -5387 12295 -5180
tri 12295 -5387 12502 -5180 nw
rect 13004 -3250 15500 -1750
tri -9464 -5889 -8962 -5387 ne
rect -8962 -5889 -7342 -5387
tri -14504 -7302 -13211 -6009 ne
rect -13211 -6593 -12382 -6009
tri -12382 -6593 -11798 -6009 sw
tri -11793 -6593 -11089 -5889 ne
rect -11089 -6593 -9671 -5889
tri -9671 -6593 -8967 -5889 sw
tri -8962 -6593 -8258 -5889 ne
rect -8258 -6593 -7342 -5889
rect -13211 -7302 -11798 -6593
tri -11798 -7302 -11089 -6593 sw
tri -11089 -7302 -10380 -6593 ne
rect -10380 -7302 -8967 -6593
tri -8967 -7302 -8258 -6593 sw
tri -8258 -7302 -7549 -6593 ne
rect -7549 -7302 -7342 -6593
tri -13211 -9424 -11089 -7302 ne
tri -11089 -8011 -10380 -7302 sw
tri -10380 -8011 -9671 -7302 ne
rect -9671 -8011 -8258 -7302
tri -8258 -8011 -7549 -7302 sw
tri -7549 -7422 -7429 -7302 ne
rect -7429 -7422 -7342 -7302
tri -7342 -7422 -5307 -5387 sw
tri 5547 -7182 7342 -5387 se
rect 7342 -6016 8835 -5387
tri 8835 -6016 9464 -5387 nw
tri 9544 -6016 10173 -5387 se
rect 10173 -6016 11666 -5387
tri 11666 -6016 12295 -5387 nw
tri 12375 -6016 13004 -5387 se
rect 13004 -6009 14504 -3250
rect 13004 -6016 13084 -6009
rect 7342 -6473 8378 -6016
tri 8378 -6473 8835 -6016 nw
tri 9087 -6473 9544 -6016 se
rect 9544 -6256 11426 -6016
tri 11426 -6256 11666 -6016 nw
tri 12255 -6136 12375 -6016 se
rect 12375 -6136 13084 -6016
tri 12135 -6256 12255 -6136 se
rect 12255 -6256 13084 -6136
rect 9544 -6473 10717 -6256
rect 7342 -6965 7886 -6473
tri 7886 -6965 8378 -6473 nw
tri 8595 -6965 9087 -6473 se
rect 9087 -6965 10717 -6473
tri 10717 -6965 11426 -6256 nw
tri 11426 -6965 12135 -6256 se
rect 12135 -6965 13084 -6256
rect 7342 -7182 7429 -6965
tri -7429 -8011 -6840 -7422 ne
rect -6840 -8011 -5307 -7422
rect -11089 -8715 -10380 -8011
tri -10380 -8715 -9676 -8011 sw
tri -9671 -8715 -8967 -8011 ne
rect -8967 -8715 -7549 -8011
tri -7549 -8715 -6845 -8011 sw
tri -6840 -8715 -6136 -8011 ne
rect -6136 -8131 -5307 -8011
tri -5307 -8131 -4598 -7422 sw
rect -6136 -8595 -4598 -8131
tri -4598 -8595 -4134 -8131 sw
rect -6136 -8715 -4134 -8595
rect -11089 -9424 -9676 -8715
tri -9676 -9424 -8967 -8715 sw
tri -8967 -9424 -8258 -8715 ne
rect -8258 -9424 -6845 -8715
tri -6845 -9424 -6136 -8715 sw
tri -6136 -9424 -5427 -8715 ne
rect -5427 -9000 -4134 -8715
tri -4134 -9000 -3729 -8595 sw
tri 3729 -9000 5547 -7182 se
rect 5547 -7422 7429 -7182
tri 7429 -7422 7886 -6965 nw
tri 8138 -7422 8595 -6965 se
rect 8595 -7422 10260 -6965
tri 10260 -7422 10717 -6965 nw
tri 10969 -7422 11426 -6965 se
rect 11426 -7422 13084 -6965
rect 5547 -8131 6720 -7422
tri 6720 -8131 7429 -7422 nw
tri 7429 -8131 8138 -7422 se
rect 8138 -8131 9551 -7422
tri 9551 -8131 10260 -7422 nw
tri 10260 -8131 10969 -7422 se
rect 10969 -7429 13084 -7422
tri 13084 -7429 14504 -6009 nw
rect 10969 -8131 12375 -7429
rect 5547 -8378 6473 -8131
tri 6473 -8378 6720 -8131 nw
tri 7182 -8378 7429 -8131 se
rect 7429 -8378 9304 -8131
tri 9304 -8378 9551 -8131 nw
tri 10013 -8378 10260 -8131 se
rect 10260 -8138 12375 -8131
tri 12375 -8138 13084 -7429 nw
rect 10260 -8378 10962 -8138
rect 5547 -9000 5851 -8378
tri 5851 -9000 6473 -8378 nw
tri 6560 -9000 7182 -8378 se
rect 7182 -9000 8595 -8378
rect -5427 -9424 5307 -9000
tri -11089 -11546 -8967 -9424 ne
tri -8967 -10133 -8258 -9424 sw
tri -8258 -10133 -7549 -9424 ne
rect -7549 -10133 -6136 -9424
tri -6136 -10133 -5427 -9424 sw
tri -5427 -10133 -4718 -9424 ne
rect -4718 -9544 5307 -9424
tri 5307 -9544 5851 -9000 nw
tri 6016 -9544 6560 -9000 se
rect 6560 -9087 8595 -9000
tri 8595 -9087 9304 -8378 nw
tri 9304 -9087 10013 -8378 se
rect 10013 -9087 10962 -8378
rect 6560 -9544 8138 -9087
tri 8138 -9544 8595 -9087 nw
tri 8847 -9544 9304 -9087 se
rect 9304 -9544 10962 -9087
rect -4718 -10133 4598 -9544
rect -8967 -10295 -8258 -10133
tri -8258 -10295 -8096 -10133 sw
tri -7549 -10295 -7387 -10133 ne
rect -7387 -10295 -5427 -10133
tri -5427 -10295 -5265 -10133 sw
tri -4718 -10295 -4556 -10133 ne
rect -4556 -10253 4598 -10133
tri 4598 -10253 5307 -9544 nw
tri 5307 -10253 6016 -9544 se
rect 6016 -10253 7429 -9544
tri 7429 -10253 8138 -9544 nw
tri 8138 -10253 8847 -9544 se
rect 8847 -9551 10962 -9544
tri 10962 -9551 12375 -8138 nw
rect 8847 -10253 9424 -9551
rect -4556 -10295 4351 -10253
rect -8967 -11004 -8096 -10295
tri -8096 -11004 -7387 -10295 sw
tri -7387 -11004 -6678 -10295 ne
rect -6678 -11004 -5265 -10295
tri -5265 -11004 -4556 -10295 sw
tri -4556 -10500 -4351 -10295 ne
rect -4351 -10500 4351 -10295
tri 4351 -10500 4598 -10253 nw
tri 5060 -10500 5307 -10253 se
rect 5307 -10500 7182 -10253
tri 7182 -10500 7429 -10253 nw
tri 8131 -10260 8138 -10253 se
rect 8138 -10260 9424 -10253
tri 7891 -10500 8131 -10260 se
rect 8131 -10500 9424 -10260
tri 4558 -11002 5060 -10500 se
rect 5060 -11002 6680 -10500
tri 6680 -11002 7182 -10500 nw
tri 7389 -11002 7891 -10500 se
rect 7891 -11002 9424 -10500
rect -8967 -11546 -7387 -11004
tri -8967 -12502 -8011 -11546 ne
rect -8011 -11633 -7387 -11546
tri -7387 -11633 -6758 -11004 sw
tri -6678 -11633 -6049 -11004 ne
rect -6049 -11633 -689 -11004
rect -8011 -12255 -6758 -11633
tri -6758 -12255 -6136 -11633 sw
tri -6049 -12255 -5427 -11633 ne
rect -5427 -12255 -689 -11633
rect -8011 -12502 -6136 -12255
tri -6136 -12502 -5889 -12255 sw
tri -5427 -12502 -5180 -12255 ne
rect -5180 -12502 -689 -12255
tri -8011 -14504 -6009 -12502 ne
rect -6009 -13004 -5889 -12502
tri -5889 -13004 -5387 -12502 sw
tri -1313 -13004 -811 -12502 ne
rect -811 -13004 -689 -12502
tri -689 -13004 1311 -11004 sw
tri 1311 -11276 1585 -11002 se
rect 1585 -11004 6678 -11002
tri 6678 -11004 6680 -11002 nw
tri 7387 -11004 7389 -11002 se
rect 7389 -11004 9424 -11002
rect 1585 -11276 6049 -11004
rect 1311 -11633 6049 -11276
tri 6049 -11633 6678 -11004 nw
tri 6758 -11633 7387 -11004 se
rect 7387 -11089 9424 -11004
tri 9424 -11089 10962 -9551 nw
rect 7387 -11633 8840 -11089
rect 1311 -12228 5454 -11633
tri 5454 -12228 6049 -11633 nw
tri 6163 -12228 6758 -11633 se
rect 6758 -11673 8840 -11633
tri 8840 -11673 9424 -11089 nw
rect 6758 -12228 7509 -11673
tri 1311 -12502 1585 -12228 ne
rect 1585 -12502 5180 -12228
tri 5180 -12502 5454 -12228 nw
tri 6009 -12382 6163 -12228 se
rect 6163 -12382 7509 -12228
tri 5889 -12502 6009 -12382 se
rect 6009 -12502 7509 -12382
tri 5387 -13004 5889 -12502 se
rect 5889 -13004 7509 -12502
tri 7509 -13004 8840 -11673 nw
rect -6009 -13278 -1783 -13004
tri -1783 -13278 -1509 -13004 sw
rect -6009 -14230 -1509 -13278
rect -6009 -14504 -1783 -14230
tri -1783 -14504 -1509 -14230 nw
tri -811 -14504 689 -13004 ne
rect 689 -14504 6009 -13004
tri 6009 -14504 7509 -13004 nw
<< properties >>
string FIXED_BBOX -14504 -14504 15500 14504
string LEFclass BLOCK
string LEFview TRUE
string gencell sky130_fd_pr__rf_test_coil1
string library sky130
string parameter m=1
string GDS_END 10392512
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_pr/gds/sky130_fd_pr.gds
string GDS_START 10385804
<< end >>
