/opt/pdk/share/pdk/sky130A/libs.ref/sky130_fd_pr/spice/sky130_fd_pr__cap_vpp_22p5x11p7_pol1m1m2m3m4m5_noshield.spice