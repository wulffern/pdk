/opt/pdk/share/pdk/sky130A/libs.tech/ngspice/sonos/end_of_life/ss.spice